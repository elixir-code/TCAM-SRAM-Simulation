`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jq4U8SYlmeDot1icrfF9XRnxVW5CPZ5UPbimy+m7utKctveEYn6XYZDaup9hluKggqOyvviBh2QE
JIr9O0IzHQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pIO5uLfyezx8Dajmav/cQG88Um/xDreFf3DYR6ey8jIWX0bzqOFMlAd0vTOsLOoohW22t30jOExF
yJLVktsoEeJup7larNrizmv/+4+7iJMW1qCVDur79Ai6snbQZkfnmj9fu+mG4fde4DPk1DgLL8dq
yXUD+sC36N7wO3B8POM=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SwYrxaOSAMTi9JzkHg2qs9AGgrExG6tBB1a1AzOTCJrIvflaOXyYfSjNfFLxRzdnP77tXQrQZnmI
gyJCOmoEtKsZyCLXG7pbGNogXBIBFAHdKn/UJkJ7DoaJM3+mcyYunHjc0m5gIUTgrmArnfkEH5ui
V6EhO7uL3qC3b7cbKas=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0jo/6ic8SdW9px7e+llh4lYUnLwhpkx0b3rNM+RWpZ3CG+W8z+YnQOIOiYHzox47dgcSCRtG0Bec
JpqXrjCWGSthcc0v0KGbt0buwgfWF6SG6+BjufYKSqLYb/+S8wM8atPSnKTKmAkx0lQ+QaX5I9ZB
DUa0CdMwnZHNZu3wN7NmrD3LlHqgqxbwtniFsZjN5W7kWN1uaamygZ8E05RFohW/aMGs+TC4f7SD
0Hd2b3O0RMoe6Cyc8UhJ2t4NZzTa1I1fWll8idRFuwXoho5U1jA3JnrITByVULLAeoUB0+KxHswQ
iih0JxSp0L2b0/oeGtl3602IrJtns579M30LtQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KFi5wdJt72ZU98Ur4+E35GHpQpBayCTw1g/W1oaX0QzRvHnwY/6jXxube5Rf6hcSB9NOGOomC7zh
v5dYPbBCF05VAvtxUSdavTAoV/BIN7LSRolqTouxUH4/nHaUBoX/Cfcr/654vee7IWYiyb4uUdKt
8Hyqa7UCe3id1xuksaPyaC7E7nsgeJerjbzjQanbtDejvbtbBqz9KJ9SwS43AvubuHgJh0xtYY4S
NbWmPB52wUcw6nd15Bdnw8WQPDGX5+F8EPp2nS9/+WVxk2BGfexs1Uir6NGK272yJZZzD5naEqLp
4TZGUDz6LHoR3U0ALz4dSnGc8sElXvplmkmmjg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gYR+foCWmz1ViISiWqotJBMvjLTbbuWjiY7ATvQeEoMUeIzunTATrUk5tTwkaU1Yx6vCdbe4osdQ
QaW8FnLD1ymJY/fdHXYi9SJA1Xd6Rwwzf/9HScMq3fg2MKb3RwRDSMpYakIg+hz8lmD6T6COR+uO
jeJedPWUqIQPLhxmMXDXIcBnwu8SikSjP0n0A+JKXUnMUDFyIX8lv41kN90e4vLcUkpiARxxw9TJ
J5XRhbG2+ynYoeBl6VYAbpATbua+zhxf6YX3MNI6QxOuzLYMAEmUS03kHXaYil7DTMxcx1CBBL3C
NS2HqYd8g/rl6NJQVl3NgJDJSZ4NY2Tker191g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99168)
`protect data_block
Pa3ssDXuqNJDTpksuMbG/Es9F9SDEUNxjTuZ62HteUyz0pAd9DsyzvmkkGdGR35AvO4Ncnf5oz4E
j1/bztFYMjfV4an4onpJDXdxHfSQHIxVa2hoWZAQhOwJdC75bwtXCtZ0Iqjnk8qCx3YYwZNNjZe7
Ck3P4q+V9w7fZNUExMK2tBHKcDHfD4KU9N/pe8MmNX29q1YQBW8AB6uym6hX6r15k6sKrCTOvVsR
+DCbfK79Cgjpy35Gx2BPJACMrvrucr6SsEsv2ojdQLdcTHm7psaLTBQA3PWtIP8O/s3hXJzXWasm
nc4u2HTWmCSMnSc8okk3BtdWLoYnzHDHJrD1bpCl5ZZsW98VCQ6ZO3I/DTONnXPNQBqE3pNv9Wjf
K3OSa0w4kzPXaeqKkjCpcvPaekMLOvxgpP0udV2jrYPLki5jwci9ooeeVA56u2yF2azZNmbUddqz
rmm+ff8UbeX1Um44SE4Sck/eQDDGDLXkU7tV0zKs/rsP6nHDUCoecVBmH5r5sXROJK2UTd5OgNcn
MNOuJf3Qd3a6TSXY/Y+ryGsMT91CN2JzGMhf7U9Ctri7SLNazZyijUsK9G1sseeAuFn1S+RHpn/4
jDXnK4DqtEeMJA1oOps/KwAjC5XqWiFSdIMCZ0Jtx6CdMcZ0S8RrXVohLICWMtpEVhX7H8Ix2sBO
UGtP5bD4E6nv5hwPHOpfbOufngb4pS104spdN7Vm2/79e1cgbiBOxRWoCo/GVctJa/4A0NBQzxi7
8bLjPokK5+APDyrnz7v57xnwkCSa2OxDTPwr8jGlHEo2sRuHCUcVHErsQapDel14jdOnkoPTH+X4
F/8WTha4NleaQZW3UxNW8DcVQMMmWvlI8sVUgEVHrPHm5EDCVyhRG+587ThYTTKYCGPQm8A9sX+a
G78RY1Wa51zoZ8iZFkNUCMySs8LWTX4WTF9uS8izpdgS4AFLbXhD6tMh3plGFXx4s9KV6SXoifIt
4/Eq57BcG/YjDyj4eClqAjKbHCFohfJZA4iRzB5aKbgtxwIlZIhUor1T5xb1KGX9c42seilFJi7I
dQLxoQRN5d5dufCI7hl0UphszcALLkMJjXzY/mE2TgNT59KHKQ6nRzsUu8UoOp4LJRdGSa5ndKSq
EUCZIfyK5Gavf9UZdeXgSGvl2DTH1vEoH88iV7e8tEtlPY0PhHHswp1/uaTyunQeKtaEfV1HWv1+
RR//3H+IOl01uKmTcrdUuF2n1shJZsLPN7ui/YNnpeKttNuq+TrBMCcHYYwyBISJhK2Xqy7TtwLZ
p4jqiRNv/ElAzL4oy/gzwg/+HxIy8/U337S+tQfaRO6J5YS5Pw1qYLIoH1L4/wcw2vGMu3y2VZpo
UNBuzIqGrC31/+EnP9lmxwT5gtRAM6DnU1USMfGRxho7+KhhsDECrDB4Pilf/c0m6lzMvf1qyD+5
pTsN7LyIyO3Kvkig1o5HHCBSiqprFKSzRF9/2o92kvjhPPvpaY7WmTNia6ZB7+kX+d56r1w3mAFp
pmAWAi5CVSH7mbsfjIwTnaJyzOqCxtfsVwtNaL3y8iLp+23i83YTTYYyYSll8AqiKWU6ob8eipwc
PMNURTu4FLOAhWCAJWeWNPJ6VRGmNtqNbk0i3qWknVcTYldJvh7XBiqzkdfuwMfxf5sxtyvQvaoA
c7tDAJ00uYMzBMGM/NqUTC/1ANLkXzdjHTV8VVpfK0qfqSETVb7HcRdcxMnPkz8Fq9+NHxxAxs+p
nU1aSKQOtBZLrywOF4nQ/3nMCL3ECMQeBtAz8kIMMO05ApCnkx3pKQxRiekUDPIFMQjhrxMCXHYG
8QT6zmd29s3yQ0j/zcBFP+UU1FxNNc2qYXRITSzKLnlgRp6n0LjLcneJQ9Caqf1KcjUrsQH6/ixD
lJvzdUT+xYD0QZpOCn31/r7yGQH66wTNkciC4a3aivus3IBpgLst788TXXR6jsiBOD5BDIH3UZXS
aNcmyGeh55e1DfX8KoVEJXsW53MjXwOhhq+oATEFMG055rREPO3kEj7HrQBWYOIpkkFRp7qlvByB
OFR8mZhjj44YLzUvIttKNOIgdC08bWQWs5I8SHnrW6r4crG9Dz3vM4iHBsLn7hiZIgvNcyWeeahf
p1Bl88NEQGCtA95PQrG/yh/yFbsZxZPn82GN+3panvhNqVtshRV+3oHrS2t0/B/KfmRkPooGVoeA
/aSt+NyYhganyhK5RtsosnHEv0siIOdh9aPBZBz/K1rJ07kUskLoTRknssEOd7gmebPkiOzI0tub
ep1tfUducNoJ7+zMJSsNZuFGHzsZKCw1M4qYXpOsAQYOMd7VupQT+0zJNIHLEcRG5q1oqfHNJgRn
wjL8h1SYC8o3k/TIglPeuRy167Be/fj4QmIQ9lsh2pV9BsNnUFU9Zrx8TBR1LRYOg/zmphhwCqj3
PuJDQzBiGGhka2/egpMa3jlZCE2xIS9dXfp9FLENrlfbrKep1mAZ2MqVwzXSZzbnW/P1sjGLAJ0q
vwxnTpn0CZ7PLkwwhZl5MfhSv8FB6svEtgvdVV42mrsusWXwq4SLUi58dMySStZopUttNlgWOgAd
pbqcmIXaVD91MswCI/chWOTYp8MMMXZ/Jt86BI7kshjD8Ck3CvCeiuKWnecPv36U+2AY0k0st5JY
V82K8p6tA3sFWgeyJNo+jen/yd2BOnnUtrDaAZC6y+IZsK9FASMJF5Zuh+fAmEzTlk0I/gjCSbg3
mg4UOCOegvUDWLi+t7FVCeC0P/Aie3+55ofgMzfMIA1Tcaoj7BZILUZod7R0PLMYa7eGfA8cauMW
2QKNuWgfh8d7ZskLyQYKazS7kNfR+bWK11S1AVUwaI4LJAFVFUg8UujVr4Czj5UGh5S7XbdngZHb
KTq5z/Og4ieoY7sFTpHrJlA92ZUHIwX3/B3E4PTI6pABuuo0jYOvrYUDX1zSU4J7uX1CJDB/i592
2ZMLNSnjObLp2tNgzHzzjgzvj6GxxWGsvrt3h6UbFonbrNe5U9Ib7sRTXKlumH4vx4E8pJDaNppZ
PLYmOl31qeFecjJw15tJR4rVI81YR6Zs3KaU/3FJxtTIH4EaxydOjFCSQ3XUYlUnUyqgixuxE9Uo
uOOlIX3QWiAVL4ta3TqCkc2dFxGRN9kD23c4mdOoAAubH67wzvILQa3oEpcofLlE+crhu43g4/7j
cnOk2DFciFKKQoj2js7D8pu90Pingn7zYR6apysGjHocSSwpMtuADpY22HC8h3wjltDiFa4WNnhy
ubriDGtyL0ygm4rhcNGEYrjlcJL3Hm06XRjwXMMHH2S04MgZmwq4dRF8piGN04Txbc+Yjj6S+TAV
D9L9FOZXxTRjh1+E4yFp0jIOgSUj3KlacObgdY/wUqDb5whYJMFqVZA1Hlcsb9SDSLfwQaCPYSiQ
Ru9EM9OuT1lDUjoQQ4XVFy2jPQmy4uaOjT2eBRv92KnnuWcf+32UD+n/Uhfvv/YD69oj3+SKqIiy
tlItU64cVhggZHI93MXnKM0tbK7vNx98jm+hTqToI+1dsco4idG5zkukt8O68Y3ZHJs5uJDJGnzN
O5keWRdYBfjrN7qk+WioUKXRlVXk3pnwbn4xFIpCwSSl2Olta4Zo3ZddRPGb03aJUspnSez1b3KH
b2qwVR2773Fxz4L9CJ6vQtyINU0CdRrxmgjoObFdfHhWYW8uYF9vVYNu9BlMjGT7zWqsvLReE30j
6AlrBL6nH/CgDkeyp7eCGcF0OZ5HI93QvL8Fq1FBp5jyOUmz3s441DHRP2dnSFx8fqCtc3GHzVjA
y1INB5RoIjNNiwij+W7sgplRI3zJiqmS0gdPwEghY0jGjTz5YavfktiWvDLKsCkgA2V2GSnXvqVN
JyYxUtKfg1TFHFbIDoW22lb9v1KNGryGBzXaInVig3A63mw5MD8sSs09+UVlBwpRi+nMlbkImQ8f
gBoCLP2qF36eHkcJz4c1zCGZ0DdckuSV6Qt/jyg4c0YjdFzhtLN4IlhmtW7l3gRinDD8NjIMiufB
y8xuMtgl6RSXQeOocJX9NOrL8ioY2diIAidJYeXEVsALSmkBCfFX9l+3zGury0LS/p2H4nTp7WUv
/cbnHkhU9Syq1nOHEdHycf+iJb4UzLZR7lm/0JlFhI1z18t+oJD5i1YT/jFrQCAjYACGgvXuBiAG
re5M+mGZ+1R47Fx/n+KdKmPSAl6XOeuKlkTjuawEPHFQe8Sp+uk4bwuVS5uAurIisydui3TL0C0f
c6q6ICUJFmnbzlGM6jhoHpXPPMLyJ0iUzJzGR6pPRjLxyZ6FpwjBcXsGY4HteRuJXg7xOykxD3D1
gy+DpbuQUovPSCELjKp/jHnW47mRGE96FIFrJlq0ntXTbrcnDX0M+OBWCDYzLOTRgQYXwqZvrkvV
rgjD7l1gNeFWDpv8srxbD470UcoMBROWX/yzHmcjDrGytyPE+0d3g4egS+i2bd+s52OzwxIIz8tt
lHLvvnBgonN2ccW5aJ16o+H4ZUcdQF8WfbaQp6R6tvMuwNFPs7uzectoiCsTu8Owg2jwQ8PQ+4HQ
USQDzMxFNlyw15vDRZFjoZh086DXxxRI4hb5bCytaz2tCdr0FMcdTydblqJ1qI21ASk4ZxU63Fau
K63nfuutMwuYD8Ci9ZGRSSjjozRp0MN334vpLzBOGn4AzV09gW3oK9r6R4UycRJzFBBB/GEgmLe6
R33wVcAtilyDcwfmPdbT7YE6X4hZ6bTFHPnd3LeJ6AzFLqnLUe+UquY/ZnlpPr3V28LFbpAgNQ3d
5ZIBp2C5Ansil2XxO5fQL7zMX6Uc0gmhFkGIJacCK9DAGAP80LDKZW5tOCZRra5meIGgs9EBnFJO
OBYNQ1oXIx66a2FU381Yh1cu9L073dJSi3lzZ8d5vdiNQop8O3WNDCLBY+e3l0Kr5XLzEF156ehq
WmHOmgdigNiKce5aa/kozt2SgOwVXV2bAoY6gW/25GgduiaS7rIsIOZscSWCSHrtjttBwdHSIRRg
5F10kooXBm+EyEbKyXWBpRMAtz/E40GcxRsapThl+giwz639UDvCmfyfi22tOe4v5HXr1Tciy9/u
rynbsgrUUoaf3z9nrf1+L5RIC9/V5nxxJX4S9hWzOwTJzCytzK+yswTXdQhD6air8GKKEYZLwQOt
iLC/twYez48EY/nHAgpJKAHZkA+umFKcTi9vCUjevDRDs+IL5PUwwG4QdQVicKnCikUrCwdeMLY9
FVjjnIjC0axrBCdcoJrDSkejYslarWskKCY3aJ1zuBKueEclOTauol/zBHiYEtetQxWF4aP4HP17
lD4veP65girfV/UGBRdHji1AZhdcuMoRN9v+OUOlazHvleyR5SYUYc8brp421nZGYzm9i0L0MuLK
bBiPVWvoAtnzysx4VAWQ/kUZ+VK1VxHN2kqm019IIsXj8GcF0PwKV6Tz9Z5d5ZE4FQlFGsNbFcEl
587iLkfastvFwf03ICyTGRlFl2KbrhyWPulaBfJcZ5yYsgTvaGjTVmDOvk9tLb8b99MxYE5EDa9e
oJGD8HAmSs7HshrSJvA9ewTO0xCRppIVyPrH2r0kMJUtW72mambuR034qz7KFdpYiAj4ZxR4vBp0
Qi0S0LRHshVg1WZWQmOmnZ3iEQL/rximtwrlSERHTg9RwdS6tNtzM2LuIpD6XQnk7fEUcyiTQ9h7
GhtoRRXUJimfyMJ1ClSZaKD5ezG+XmZOalmGyInLdK9P6yybNNye6b8laFFZToahc71SfLDQMXq2
0EPhOrtLNCge2kPUedwEmDU9EqZum70J3hSUeQwzwad/k3AjoDlt58c9kIZl/ltujNiRVIvQiZxW
shZYEFKKYN+hgE+6rJFtMHLblJUy1WTuSoy8tWNpajfxis8tp9hYpDAN4q7x4TBLEQzyFb4NUwK7
XSanVjRB7sxDAg2fCIbbsTCWT15BNsUYT0dN/H/ctuJw4EIMHWymhIBAryWQNYORCFrhW+AS6c+x
E01G/Vt3Rw3BRFcXxp36fDhOQ5JBe3oQLi8mopSbOqdLcdH0l5S+70KpK3aeAwXj2BQMCNR73b/I
fHxewgZun1zkPOFjG+o0DEn2bpFZC5+5WgdlPadiY+Ji9EMtQ8K/YtG7mg5CnHZWbgLrikw8nGh2
whKYpZLydKOG/WaJRScrTdgbIUYAniFfrd5Y8TsMarlXddx04g5/4sPwQiXbEPtHbete4BXEoPkS
eGURtXevQF9Z++61NdSab7LMS6Y5UyubGzHFUc4Pe+5+f0XUiZLf/eo2fqLxfUpbeXraGXSnIbCq
YXN22k/Or2IfRO8uC2W7dyfvv9bCEU88he2tkaC6Ez07Bpj4wQokJzNPQ5vG5BCIX1rXb/at3t6p
4ydA98LYwo3gEhjAapsw75KdH81xOiDtTLakdTKrL/+OMwGg6ZJYF0U3Gfn4FIFpCgw1Tn7wVm3c
pAkg6L+uNofXDsxNSjP3JC52ORsVMuTR4Yf8l/RriuFJyBWPo8HhVkq6JbisqfYguFauAvJK581W
ws1KC6CYjoi0kpJjnin49xR0OiIyUmHWGV+HjM03mcUp1edwNxTbROWNiEN8/Qi60ASDf1z89AiP
TdxR7X8DCK4S6YCcjhbatCXs3t7fFzB7YayY6RbntUe/PvsHYhsobcU0AN8AHZcO7ATXcUecCNHQ
pZJSZCUQdsg0CQbKGo6PvN7E2pW7ufbceqXmkqAfAvWXz0ILVwtrX8BhWQQYszpeOJg5psMSFNcT
K6yBIRImmHKq2Pp4UGrsef6jzws6xOJHg7d8rWpWqJ6SgAWv5/tSGMEZVpLGsfuGRhb/I/kk9Xbo
CxtUnDGgwXGwl3OCimay5Z53sO0ef/yLF73ZwkoQf4Q6Qhk417ErwjekIqNOAD5BHxe4j9QZ9djW
YEK75k+o7hY2UThJJLJp65U9gR1AeTyhXquEOhCn8Np/SmUq335dYnmQWS02ypC78hdeEDkaP7ok
oasZLCgiQtU15Ckenf31E1tc4An5nMhcEmpqr2yJB5JLIdTomyaglwlZoXVw6qxHMNSIKLke4x9P
WxDlOzlYiCZj432BrWpNZgjnrcn7/HMWHMpUOQAHgYoYFpXerFloR3rFG9s762zRhpQd1qO4/GGE
24tewkRxe8sOEahXMUeeAFSkgtU5M8ACNqSbavYP6sGX2dbo4BBUCxp30sp7c6xPpVjw8UT99N0/
YviycCvrBcFSEvTekrI+h/7SgPSYihIAXwq/p8wlfvb0W1V2DFOSHLxOiLVTTlSVqvJtoZWrNJC1
e32c1eMj35p08DzRAaIiRf2wiXjWM9l4eVoAOB1V/e0p+GgvrnHd6jRAMw61QzFF9u4ZfBfK3Kqt
pBCxN3VEgnBCzQsDTdJQCGThXKnlNdFr/Lld67yXv4iaO0shhyVbcKxZ1saPdAymgja1a1G6ir6i
Coq/RKM/pqcr6+V4Cr6OqfU7CGzax9qbrBJBM9xoPSFvkZWL8StNEmQnwdFh8mR1HNwik08vvoeD
Bzn43+CK14aO7+tSryIl6ZsX4uNEvxxGj7c+IcGU7+0vNYvOGC3yqVyh90ZJU6of5YkQtrCHPWpU
VG4k62qoxHdeuspJDdvJCdyavyeLY37z2cuXDXDIBeNKbEZbzrYnkwazc4iD3Hy5xKUXnsTHKCbu
FWkI/GkB6Hsh5+Ck6qOLAUY3P2VVIri4JNE9til/8mAKOBxKLeUH0V+JXQnX817h+SPKdu7/p/+k
lFctQ2XylvD1d5Ny8mQPgLfsxk+GiTNz1hfl1nZxtJ/nb+AO5qSJpSx48nsWbWK/tmQ8Hyz0C98T
4HiQw/KK3dyUEo1SldUDfrqJMsckiRaI2vw4CKBhpo5197DEHM8YECMyHk3V9HTQClkOE5bcuDY4
y3EGDJZgpIWyiycYRqUcgB3k+k4mpTdnF4SZ8+xPQpjMFcIG84XfP3AVJOvmrt8z8a01W1OdOjd1
cV7FB3iFygJvZPl+iwLyFoHLywK2pKFTJJeJ8WfwoJeqLChWWHLNBmhBXxYe9hxG58H/oiFIPa+1
X3vs5z1xjVYkGZ6DnQYL6dhqiVDmyAQ73h4tfi6yXoDy354pr+EBIqCSdEHkE0ueog+dZ0iQoj0A
yV6KCLqtYJsRAtUwkWmGyN3GR+BWYjFgdXpcXf+epIGYJ1jofS4Eoq9LEE5W9I4cbXED7wN0JFKc
HGdx3IGwkytzAVwI392V/F6jPeVRrkR5yu/SRalOiI1toNw1ItDwlvP1SUHr1cK5nAhWZ/ZmoVYD
dYyv+/DdO24wKy46AjsI9ChT0B9VueCLnkFq4a7lNhvT92HIEiZWqQy+Au1XO/dQAKy2JZkfcQ5N
hV4cGF05+mxaHzRYt7vvon7OcUTDhNBbg/puSxNOZAGPkZiko73Jc66S14HS7ONhCx+uaVXo+4Bg
nHAYjhJ8LB3nt1cov6CYGgiFNtMaepIZ4PwhY7YWgy3Hc+socQEXR67Jhkfi/QccIbG3Ly1kvEdu
XPGERxZw1mqYbAmJT9gcFOCMgnRZVpdJzDJHGSdWGfCofrNtZsToM7EZJAAmEXyyXE8R5FlaST9L
iDs0uTmoB5wGlwpom/7XUIxUurw+oO1u1aqW+cpz433j+We/6EqBnLmZXYXNzaVhyZ0Yjdq3P86N
IycUuS/LtU/S5V5HeeAh/7UaaEQs8TzQWVlmXI79oVm/FFJYqd7dLzYRN4XMdu3KztzG92vq4G+T
a7cobAxTQz7A8ThCOi6FGvp6a3AIq6py9Hdy2+1jW1jUFV7LOEeD3GVJai4dUZuO0LlzPZM2t4Ls
zx/rGh7QVbJI8vnhi0iMsreJzj/Vwjci2GA2whulS0UT+WPgUMRda9kzScKoZPmB7Yg2zaTQtBKn
h2W0xcrjVWCpept2sGEG4qRlid2XpvUfek22K8hAddg2Oi7zKEwNU24iwvICsgcM8n9ZON64fIeC
YMIy8VL55W2MV+h3XFzGs4N24F/Y6xSIQdZim6QHujN+nhfUkL4TL7xYHwf06yAxMZrFRqYnl29v
nkQr0ji5idUpdr7dV+XHJM+F15YhsP2iwTV3tdQJeHhQ9/erTE+PWq6MGAQa+IZOKOBPXYDn9c+F
YKODnwyfV56mkxhD7nlPuFwBb5rAsyAlLB1SegbCRzaG0N7s2rIG0y7iJAqO2675V3U1s3sRj06m
/Gw5+7f/ngOOuTIyvyo29onsCSRr0bWjl6aV49fkuijox15ormY3RRIfvtvMH+nyeO0jYVKhNiXq
CbEsqQ52XWc2Tol+NQXv11hzBZo9bO/fcmHt+frI5tFNfDWbjpebr36StPHfO7XltapC+R+v/DU2
Sefff28EGwoUl6oKNs23FasaBA5bDcPbdUz6lihD6WZbYG/aW4LKxajpEJVZ//1xrN6bcZRyd23B
PYAJMbi4rHG38FT9i4SQqYRTcRSKQCqeMhSBngu8SZGus+/+W4LW0JaCt8EgrWTdQBmkJ3rBOAcG
8M9ode6oJNkPwfTIZtwF25dZvdQk9lFoe6OoyCmnBqprLuPJUY+RBpfZHn9XVZCQDBRd4aAcYKcC
ikp4SGAeSbT30zlBwh7MP+HIHSnQG5OMEBTfPcfZVMX9k7TMIILfAXvTOk2tVTtQ+eP16PGrv0+R
sgy8xXe6IYweX90d1irK/doKz2sNpQC4bA3hYdcWVkKFn9XEa8sFF7ytCvYzxQO2sxmcnCZOnRpn
xjD1A+/q/17nSKdo9RI5VlBF81VEI1mt2cIwqOz6lUmytZPVD3eui6qhvqAWY1qImp6zvQ2/W/KM
gEpndCLDyph/P92PCuvZ+pl14YOFTkm3VSNJ/xj0i3DEElf9ZSuGKHid5tDHUgttb9l6MoiGSNGA
Fkkh9YI0kQmXmGO0hHzy157v5a5is74dJiru/hOUwUOxNMNklnZm01RA/JhimUyopI4SkasbLviY
Qk12POQS9uaoII+bC/HIxZQaiRV3i22GTrQwS5sVDz/OUaLNR0rssS9ut3jzdAvW5BRJtNY6axXP
qGL/buBwbsyk7I71/vMQ8JAXGNUoLZo175nvQVpKlaWiU2165KBG/A9oK0dcBRKOsdPsM+k3nUev
dyCa204LUqZm6bdXncA1FjQR5xHeHBIHt4InbJWKUjuySB1nU1oI9qRuvSuxOXsvS0CBGuPTtj53
v//OEAYx+9Av1DqeyFrH6hze8pKprCfmjr2x0g56wRZU3UbjTIm5G0/WC+sgwaTVmd+0LjrxpAwv
HLPAqTTGFLHC6nVZjEnnPLh+wiEuf6ancrNyMlh++kW/r2Mg8WZEAxBz7nniAzM0bLmZqSOIi5hF
M0AGSspgy4t9y/E7Xlus46nDx0+ZBqg0DZk7i6T3AsfYAJlRmBxlodZOc/RRxPPzqe/kZr8CHkFu
WsrE4ZcPXWxxTNAuvcwlPwLdRSu8/LWYzukiOxFGKmoaxRwakOxR4zWjQFIpyc0vR9I7loxamR0b
JNVqG1mNoh/6OGAfgpzRtZ9gpdKY4+TzIs9w33EFTRjQevzXxG0KKxu6fQPVwv5mbn2ke+k3bWX5
0MWOlwP+MZQK4V1rJYVzXo2f8ina7rIbDWgvtYX7jAtEjuWFxPHufzJhnMqIVTK5iPB/yJYcUpY8
96deyw3Q+NeU2BUfkoyIXPHfoL5OvgLFOAKI0y6lMCYJIp3qCLc0rC+/2I8Tj/IIXG0V3Car1CEB
mgBevqjFAf+8+vWtbVU+4lHP7xh5gdKNzrOle15ypN1NFH6R4duzA6CbcyD0S0OLkrFgbqU01iK5
OG7KVYTgHLjMjRTkXrzZC/UiBXiIECAeIhh7pLkORpm4ZFnCKQowZ/wmepyZdG1y0zbVdQ7YaI1w
rmpHDegOUB3RTCW0XaWj7BZeWlHNk+gQtjDyEBlvXW6qjFsD5lPMODDVqI72Be+Jtw/+G7tHPs1J
APm+T/umoh7w2cLuvbGdD3JXh61T/mWmW9GGCiM2VzGPQ1tCnsixeLaOrutFAZcxeQdwjWGCML4n
MGR2gBLBoYykOVoHrY48LpRQqI8Imje39DFyRaefN1CR61jorSOuf3Hz5ORl+Q0ynEzhVS0ANIM6
JQJJNYUE5EsonAq3ACH/AjZdYobSCef5Yh4xmFGE9A2exnK56ponWZRJQtaP3cCPW8yuF7Fk9rlB
1aPgx1mzHQ1r7xjYWrsz0qCFxeqUxHyW/LFj8JjuDIWOyrndK7Yi2WAnA3h86DtD7xhZcEG7U148
jsi5r59GIEefCxm6kcjR8bDkxu3Ng8/ho+cNIoP8mOQ0N3EaUCQRNcIoxxE5yvLPvW66LuUJJII9
/OhorMhug1w3BVF4skooDNUrPwS7wZQl2AGMJL5FXQgCs1KxF+dXP0qqBXQkSoc0siZvzi2CE/vK
bIvRZ66DC19i/dAoRWjSPJVad5iy5y/C8FUO3bslq3XoyPoIXZVTEA85LgGb1ryqZPUpeplyAzct
VqIs3GXrD5lZrFsNQvq/rRGGgzuOwFcOohdYofnBZFO6hOHee/HdJSFpObC0zKaE04fHNo/9hGk4
rQ0iAJfaQBvc1ZILPIFSUbhGMQXIPAK9TwD5xep4ZV2xj+geqUEfGLtIY9KhkyPtBsH2CweA9B6f
RboydZBqIT6fg/JOa0ZZs5exDhVQjDvonKRwwbUO4WQTIu4HpTxGqCv09lQXMEMlU0ilYkmI//Pv
Ostkdqlu/N+k233YscJksSB3qiAodpeDex5vc86DXd/Cr0z5mmN0pLnA2SU8U6+ZTZOMfgM65fVi
OPWoOeImZgr6vfzgVQsrdwe6uj3dggnIvhbNVUa/qTPDe/Ixwa9kshFQi9uWpej+El1lIH2R7Pu0
0RdiOFql3B/tuXfjz4qjMqTx0CLfcplbdG2o2ajPVj44vUjPvlABZfgnRQWY0r+kjduQqY6S2UjO
uhDGK+CE6PMBfIZLu2TQlunDZX2IFV0DTUo2kelAfoYDzXqhcBp/b3LpkWju6QQ4nAQmXZtuHXG/
cShlFGTjzzUGtTdMfcuUJg4Df0Ua+wlRRvgEZvabUOJiuE98aI2XLHeso9CBK+xin6dZKHHmoB/r
XMQ9fGsPq4jYB6QmHi/YLpsxU9TZRtddqLroRXm1h79p92oFBhA8fDn1yoyAyvO+Ne1aqTdwFaAH
CyPykaOfSmpzHkZISoX0/946cXCaK1liCZnGXQLsF8qVdXrLHA9EkK2ki5D1qY+m28XW6QCl5sgT
a1oWyPS6czA27KsfObA2mPz2EswKjcKodvtqn2a00jGbwfqXGugJ5JWs172I/7abTMIUUyLAg2eZ
tSACw6bdYm8VJWNmZJraXY0PcMliETOroor1xGHOKUCNRtCrarrAwoGl8f756J6awq4wCBEJwdO5
UiaojusRPN8Ic4sBH4hEKihVbOP6Lk8cfh2FejNlvCNYQw52/qFmy35mSf9n62r7HKh7PqHTIuRo
HXRSa9kaic2AbCSScGmpXkrQ48ZhAR3/ooYThn/k089zE0kUIOt5BWeUs3GNz3TTlwX9jLBeddOO
Qq8PS3SZEKgr2svjEhNhGKANDSELs80CErqA7bXYz3E+WanKJQ80pqGcnCk8I2Ni4bDSAEGAna83
ZPJZVLnu+zJ2wL7PqU9NfLPdPVG4P6tj1mghwhYxq9DNCbhIgD7edqmZCTYQ+9Pzj9reVRU/qt9A
+MQ7CyjWkCtTHNXPtdN3cWdfKYx+iqGGHKy7d/eW6lr+9/0sHaLFefploG9O4CX1T6RDJCmasWAZ
ySUSDOVR8a0+lnGCJfUogFJd4R4dcZMdsysEVdrE3KToImspBHNSa4Qa7gn+qzLNlSC1p9b/qKsO
5dEn1KHSEu1zXYHw7jflKXjmVaoibjWbfixaklBYZde2cwzU1zxIZflJUHz58l8WUQLfFoNxxjFr
dp2wh0p6erSMOAOyBznxUIpZlldr92PQXdn4qaPIrfxSnU79CJoWgUXFMwAorX1r5ZMwh0ad66Ms
3SMqpgtMHk17b6sTCg71fJgmfKA/uZOJdCDLwqUtfFNQh2pIp/hOJOit8ocD/1lolJ1j75BoPCYY
t6Fha9dCIncw7IOjRAmU6NB2+sD9bd24yFp+XJ7Da3801xHXK0BR9zbh1VpcjOhSZ1avAHSq2bU9
iepvsLHp7Tz4km6gn6jcgvF9LLxUmt3yV04VCWtSKsMsJQINqRI2OhU08AOYGmMJQ2P9kE3BMXr6
DLyPxCApY6xuSY4KmxUR7jrZhPryvjU4mWVHw2knBM5XmyiG3IUpWo+3ZWHGnL4AFhSfc2y+l/50
eSN45jClIQoNSzkbdcQGrVa2zG0geXEmlEr/ovW0FIADuElyByOl814b2LyDUV70f5O4OBD5Hbgk
mYmwBU/d3suzp0iwo7KMnx6ciJbPeDFW0kgGFyJN9++G2gyjjQZbwAogZemgsgBeD2MO9pqPHzwP
MSpJPSf2pn2PpzPPWLHkNz7borG84aBaCUUbSskdJ5v493PsbDGrfdI3PnSKq9hJ9ZC2b+rAGfPE
rEzZiMVis41T/c/uRIpHaHEJsQaYfXjJ02Ii9PFxEKlygw5wOp3zrog3AXDBEGuja+zn0dWtfuwP
EMTB7mNLe93jwG0Xms3ChKx3jgy0oky/MdaE0iMNVq7j4f2aoYlW4KFVR49Wf0eP52D1v/zKckua
s9eAiWE4Wb3I9Tx3uTb0pDBH+yEm7j+PxzQwyYFjorJbuAg2IEKvFIBTHsVn+yeBJs3XMIvJSdaX
3UqaIGmlESGKDUfh/Yxcl2+9GBOIQTZJVuHo6Bwvw+ao+t6H4eC/s8jkEEWwDvzmOLw2/hSIG+J9
Y5x9eKnlB2R3lHkl2kyyet0ty5LlHV8t44Ad5t/km33n+qrVwxwY0TvSkF2IVkPgIAkJ9eJ7GLZN
x/WKgaqXGL3uLzJ6wpmJZdbXoUdlXg3Z+FJUCySiCjoSd1W7JIKcU226QVIS5YTKtv7bO0BlxTvr
EUNXUvSApyajEaYcfa/2Eukl79H10tx25V0B8r3vkCVxCU5/5+N7GtMZmwnWzUTGwhxqIBkctHNe
3cBIefsziyA0EdBlW6nyk9w6dWpTKU+LnloaIckbLMfq+H4NAtqe6aO9Gy0xhrcQlMyYhJhcO9vz
MSGiwNICxRh5hB/toSKzuuGb7/rj2FS/zrnYsR2tgKpnnyf7AAKTXFkZomqAVEKZ0AWezzY6X4nr
113ZsZKaHN6po9H/TkdHUueAcHx43z4JIb32bkQ1cY4M+MZO2+/pdh+MEh7h4yU5QXriSetah9cr
SGmbDN7aRpd690FPy/MTKpzfLHYxOx+Qsa0Mr5t1odTztVUorrQY/GcKUdYdTycbO96tB5GBSc7v
2w5xUFHEfA1VEKcIjQohjLQo4uMWi264MpPN+KMRolPB9y6v1sl5FQNfFCIi7S9hYuOR+X+SuSwZ
IkYaq17rRDZPJgxluwfqlPNIQprxceyqpuVTeAzDfnyxuHGxgXcMDQjTkWH8fCW29h7TaY7kg2Ap
P4PNHWy7Jh8ceaaxZ6dAnElW6yW++89r9m8BGESN03f3m8g+vYhnHKxWtjr1C82n4NJRm4CHZ/F/
56Aqsi0G5S9+kvjp7N8Dt5tTnJL99RPsdEOz1lAhTUbZ1vag9/C28iQpgfltB0TA+OWUiQHquuEX
m3tEfMS2EQFHH25P6MCP37JKhzwhRFeGjgOR/ownXo7Wcz/LUP2VKTZBtSzMLuWqNKTEczdi2Ijx
kYDTu9JeJZODj6EWglRvyzLnNCJ0yBBMf3IKM4czx9VFJWqsSj6zw8qU3f8palj+OY9Yl6ZJikhq
OowvDYh0vA/eI+zrJpk+2hi7c062lWAxmq8m73ENWm8Q39M+OVK6k+tURu4nKEoAsc+A/sYgMMou
1Je9ojYEyTkXAsBZGLQwvE+554UlBFqbexdaIR0S7PjQLig/atCz5wQ5bhrZwd1fz+v/frqRsoyo
eqQau52SIr64UPP+0Sb0C1tcGf8QMUJhqPDRgzyFO8ENn40dURfMha3Q1zAoVHXMBYHAECBXEh2X
lPK/LlqpoEwNPJdb2DaJTgDuXW2v89TZh1p3+zixcmXWRDJm4AVi/n1ry4aSzFbrrUqT+K+gZT3u
zCubkpENTqMKxsodRsP3IwCLLx82ZDEPwY7u+y6HLaOt9iLwWuKd6mFKciGCbq/B55NqbwOPeYrg
ftq/B5dnRvVwlinD3MhiBNBFM4uoimHpltg6oC9hBHjnZkh66ge3yIernTc5SrlVkE/DIz0J/iqB
8kI20C1CeQwfKF+pJB9lqDEFW1rYd90m4HmkfkPsn71XK6EgDcEz8Ile2eK5FC31x/v5MhWJQt0A
rapa65jFCdEDovELkFlSJN25EM3JOz4g2ie3QRMIPmFShIakVUXPkQ047knFF88MvSlBbQHqt/Gm
ux4FGKRVq4lsneVA4t+GgYrH0icDeNo9rH1Op1REeKLNofdlbcobEGncryaDiXofktCCrF4r72WA
6hbRmdkq3qpYG7YkwStaZ0gBVcyn6RoigsRw3relaYzV4I/iciku1UalaedwLLPhP3mJHWVRAIFv
m1PvjFM0Ls9s64qlXM/2Ocl3M99ngeuHbN0tMrUC3pTaMo6oJzUHQKrGGncdxQ8erA4L7Z7m2x0M
C0J0Fw27OtT5SxfhXT2ZUCHJcdY7TUQtOuOP0y9mpwekaKX8YtshOzzHNCD8AijB1cPqn//ly/jD
r7d9SEPM5I12540d4W3R4f9oaLTDJkmrN0NnENJQ5LetnRAAhsRjXNPz5SFm1cmkfJY0rJhAlEeZ
QKQ59d1d8a82Ak5xYtj0deYmCaEcoRC/51oL3oFOkOCmsESSAprJwIbyeYdFpkYJdVSa9HpJKLGh
8mOIh4d4SiCTGqDWImoSo/uGkUMVjBBdahdXY40A6E4P6iQ6456uSoGjKCzAcvNyBV6k3Xra+sfh
wudi2pCnUQp8ke5/eJSeMk0T9PDq7NZ4ldE2S8FVtQBI+Fyzp+O4ZLjlJo790/UGDGcR4QzroQb7
i0ooz+K0BAVUnVwA6a+EPQww/hussaZzsvZxGphMG8dxrPtq5SmuT59+34iyqIYQtGvy9TAIiMQn
uQ27oVmZBmOdYI6mFAygIpSWr3ORrbDRQfuBdJUN27bdjzyz6tBgvmYlSfWhulCvyt4T8FKTYM2R
2lxOjmAkW9gNRjDXm2EWfsv8yxCUxQJ5aY1qheRzrCIpeNzJlSflQP2FDuQf6PvdfwXR/hSRYpnA
+b2q2tM7bG9wsMo/58Dg0xVgkJXI2Nu+//lgeeXOHxugNj/+mAMmfA9N+ZIBd7YzYwgMDm5IX8S8
FBaTIcnjwQTz/lrhLbnuhqXFtjxSE5ZofRXGc9n7Z+7wsGARk8ezrV3rEPO193sEOqHzjWZVvdT9
O5XOivT0oFr59sVjq0WyhEVUVmQsSu5EeaniyRu+FNOlKeQUo1/l7/3hesDmpPUQNq5/+2ndSnVA
6UDoOpo5K+be0ZiD7fLVPGFcBmZxdMthhmqsPIQrZg46+9d5kOfwkq1pEzAOMlu0v8NCNX80yMpI
MHn0NSU8qxFpxk1Y0wSxpTbgdZWPLr7KpOIB73j92/paHu5fJN0Q+xqe92Fji91WjLl1lOPCZ9mU
L3tJMlpMrVGWccx2NnaIMWBWBUA1z/yQ+3tbdoh70zGyJVIpcyPpfvyB/GkRn/pwPnNsDQyolptc
ixk7rkkN/puDlwyRgjHW6f/l47QepRqcKeoxW/wUCeJprQLACc7I5FxJBIhXNnyk5Z5MnbXvJnUN
VKH9lVzS3kYkLjXrYTbNxqDrVySiTo0ZGUgWaIge9oVbyIS7RNG8fm3Sx5B1sEXqmdCvLQCE1ZVb
NK0d1c4iRJX0iywmg0KcWAacIbOdZQiG8oc24PW1151gntqjrTFHiPLaPxVXSn+LVKWMEAPyOTYd
PG0M9t1agBiFSJsf2uRlLKiVnBVWhATMl9liMC1yx1r8VnESKEDCb0Xe3PA/r7LyNE7yfVZ1lj8V
AWa+4DscjzThxFqzA7erdZTaD0b25xGf5y+OieqMiUwZSYjOCoOy5ghpSRCs7WhroND136Jm+OM3
d3by+EuHorIxMTy+ORzDWQkWcgOwlqpPbXxkcQW7Zeqm7rVqxAqZ8h8Gk0ZteTqJvuUWtZUlb3nI
TJIiBOl/svIkZWmpNXZvjX/rt1dPwOs+fVZNsKDImdrMH12Yn1Nwkm7d3bio3P0G5fEGq6rQzKhq
eKOuv+pBv1v1myqVokwWwUrJAaitsx8Xjm3tpkUrm1yQTg5Y+CvuTP6ASphU00vQNG6CChbzaKIJ
/XTFEFbCVAV2VOA0qO8b/1735Yyqw1D9mceOjt6BX6LdRlNPu9OaeIK2TCCmgZk3NbMz3czcsxrL
JI53gAqnu+lkEKXP0AGy+F0G8mNnQFRx9tq6MTDhVMgfhUUGLwvHvC02CmIHun2CfPbXDrPILtJZ
OjiHJQMuSHuP67ZsXy+P+Nuwef6nMdsL2dCbpp4awLGt/Uf/D+8KTrHxFX2sMN8j+bAM4Se3JllN
Hshs20+nPpGzI7NBA65NrBMNcOJ0vdwetklL+14GmvtWAM+ZpSs9y2H1w4KiiEtWAlpmBeq9O8IG
/2cIiDJdbNE8F8afFA8E6lP+pe5M5VuAmW3zaVdZeHlGUS8z850lOY5gQS7Qyr7sP3Y1+DG3oqzW
Vi/0jW5C0LAvuBqKKKsOdHIlYqm8Dzq383LKmYmmp7VxC39awNQCMLBGqjy00dfFke5q4KKx7dpr
wrH/F1As3fCogCkpuj+TY38AeWre8qSWpS9vRg7DjIi7WFZPilDNDvgYrbjambHfyZEuK0Y/PF29
XO9Att8cMOz+ggxDUXfIOe12CYjPIGfr9XrIk1Hc4MZh2xZOsXCPIkRptRfSnwB/6QjZAAYYBdTS
4gWB8eFrAy8Fr7zW85g/33mSmaboJoVqEvFu8nOhDvjlzcX/WmX6R/IDkY5LcmtzY9qNkzS2CZg5
MN2QqwSWsrQFTjG2cjWXPb3pSSxZ/weQKBacfR/eVY3coLdwjG5Dy1jiXqN7zaL3J6JZmcQa2a70
XenQn8EHklAS0HbW6cnUNQSP/8XYHXuHBu8hklWgXcVuTMHT+lcwc07AWD3vNBncQfUbY7pVRsSt
n0F6Bs+/V48xtZyoZ6hgPo7EhMnDI5W0wIUjsTr3jGKB28+6u1JDAsAuSwPcSYlK3WirOA9tNZ2U
qUiQMyTnrGk9ZdJngHyOhy5GQ3K3lN6L2NX1WimiWYRxu/gGtg1itgacfNLsTETHW2uxOOlzrpwg
46/uS6TAKHKWT5drRQwq8/kX48Tg/q1Lqjd9jfrIqNqEvjvbrFBNgeIy4CkDmUOaMS2pRsSUdGtj
3zRRd7eImB8eYO857lr6hbezkApA4hAC65gyxURlKc1uW1Zx/2ARCc8jVXtCQY9Rry+WJNXw+6xJ
8aJChn+SirZXLSnf70c89jyXbOB707qqv7E2hjjySCmqsCFS2FmzJktssUj3tjk2EHRusAqcxMhv
rHx2k+l4DA3GRaCgG1U0MxQRudyowqEkxPHp8nUeqwk4DHz9cC4GVA2HWSmL/6sPYAH38zvvJto0
ruSsq0Tl8RCO3quYDtDe4jks/qimFq+62WjZdtEoqcV0oYp9/DO5W57bVadD0dxKh5FvWncPT3Rs
BUrPFFLYIYB8OjEcvlaA/u/8mpEGiojHNBM0qKSc4TJwKVHONimyNKEpc51bBA2wt5LkSu0hM3r9
xvaABo6KEUIxMZplOEmr/hnGH0qzsJmiUWBMbE/J9b7JRx3Ff4W4YpD2ZZSyRLwMry0zIVN1G0JT
PvD941C0zh9d6g8ZNWoB+riA7QTvxNSfHuwMMk1u+YxeYjXYfmsgagpZ7VfBGGkAZPq6utgSH0pT
M/dQAhGyGjsKdMTFFrm33v610OUbizESPzNhKyPQojexn0iF47kW4HWNhIFk/vhUMZML+KLp2OYO
Xrn+dsbp4UI9RsZQPkBdKJONRwG5mbE7kZLdCZx+OpiEstxMwBcallb9HNTosY1iY7nNycUlkKFp
FN8eY0RUMg/kXpFJBTzoRojc4myTvNNsH7Gexv24mRZDBNmIkTjX+03AvaoltmwKb7yE2G3oaWO0
qJv6O1Vh4nybyD+FufKuL6feQFLVFHxNa2Hh+7IeVZXVPfSCvmgf8N3H2VcPSbC1IblqsaImxKkA
Bmv5BMg7G4P11KXGODh2MZsIqfCG/EgOxqul97WAunjrVHOdkfI7ob7Cn0XzDNU7AzjxteIHzZQw
l68nZSxexMfPxWldePvhtu+L6tXDMPahWUCNYRRJXxVPOxG4mD9Ho8S6AeDVNWSseq741KbH7NGd
yil6wpzeV85aDbum4bIfoGBLe0wMgOFtIeMMgVSaQsgG3GB6ouPoZtD0b4Cbp3BKQN/ecTv++I58
dd6/vezsUthq5RF07IHvd8WfOcDeQOYzRWROjhac0C0WmYDYwNqB5KJ+jupItk6cfvucvCg/rsCK
9PYytaGJnPyjwfXvvQUVj7hWi8ztr706PkVNLEPcK/y8lAgSqfj2FRZr3vNogljEY/wDxQoaXi+Y
KA3+xCyfz6sTqlgEUe5EZHMfBXmqka9iJc91hrBZWBhbyIqZbpsk1ZZA/sRUIlcdSdO7apKAuZSU
1LZYg/0Qn5JnX9U2gd4A8RorQ2uFJOqbzLwTk1J2TWhIW9bc32349x6xFOyKiJ5qS87BNfchIZio
JUQEnszYcVUC93DyfT54W7ipb3Zezaojb2BLFoZbJD4Ajw9x1SL1i2tckUh/sL02eYmMmDfkUmam
nFifl8Sps5d49FtpFV7vv1bJzG+NyIkmqI2thrSke5e/6YhK7hHI341+/eb/Rg5GNAZq2ffWopcI
K5RiESz4Hrd7mFy55yAkXfmIDBLtVYmQITcFnhhO6jO5Ivgg/cx1GcQbTEsMXIc4bbQntnvj3jvY
FBu8lsuEp9eqZixqODWluOJg2eN5JO2Uh/coPDThponpHsR+H5APsN5xuF8aLLodz+fKL/G8zDCb
dtwVUPcUo5WkOROSxyWwXoX9Nl1wwQQxGFbd1NhhXu3aXEU/OopULD/mkJxmGdgq+bClxkQyJAvi
N1l6Yz0eSfQL28Y4aMZ7Y77EYy1fJ7B3ntnhgY/9LBZqBuAYlZDH8i3WijdMUY+pFICfLZ1e0rrG
Ugap8WZv9tBP2n/sD1b0LjjxOWq+ahMpD7pX5pGpdBUKIluVn44hEPqONt3jRtsX/+ZwBHyuB3Zz
jnOgnoAihSdDolNV36BGATGYGkZm2g9AymPMKFfATVVgCr8OuipWL6NOCxRYkNFhekffvP2vNPs5
MC/wEftO2BzzKw1Tp0A7v3J9s80z60VVurdUxiRRb/PX1YFp21ysX1V6U2XMvMXAw66pBhBh7J28
7ILvlsrzyBKQXz/8AKgafjt6gQb2IM/oadvshw0DBqnWjaHqqVm5movk8cpbP3eU1qKx5SW/QTR1
7W2cPwGmgFEShxY1OJGCQt/4eGMaDkN69IdlyduXoBjJIM9a4vI2CtBvOz5SS4IOvaSrDL/nOyFd
8WodDmfB5qOYA0YVApZ1a8l4Dki/EPbuiiMCiuFFI8/1+WEsJQ0Okt4KISUARBbFRdjXKaMuA5Bp
NP6cmhlBpc6cKF+VKHq9nutJvGGyHvJ0RPYZhunOsp7sOtbYJ7KPe80+7spmPb8YoxsBSHtHIm/f
Bc6a2tsQNKdQfvVggB9L7imzsVjfp1O24N4MVR15qmx634S3x74GAYfo+CfQ9EgmMeaNWIrwKPqv
0I6QHbrIyzFFLpVrXyRUFOEdUfXX/t9hZE483Ac/THDItT/UCHtWk9w28O52lpZz9rlS0mbFZS0i
t60rjitrvQZmDSoCgVLJxrogMhErJ5ZVyUaAZVQ4/gOE0d6JIF2u3lanu8I+J3P1A+n8fXbn89H/
C7N5+1L2RdVWn8nQdeuSL5N/gY9uYPMz/v5e2lQ7Lbe40lX8uZX5HK+YQuS1C+Pzuz8f+TOk5KwT
NgV+7+yApkOzM+xMiOCOhvjhj77lsakkOWrGV59uF3ZWaJoDNKxWpaHduNIGjQUe8/857UsvJSb9
JwjxflhH5tOdr64MSVgyxm6ocNsrkaNDIl2jSfAhBenDExw33mWt5/+49uosocgo8gkmFGsb6Smc
lbEByurfH8ZpQCCE9M2kgUDZ1wYrWUbKBPixAJMbVUsv2VsRL+HjUdBAQidiRBI5DW0pPA6/WVFN
HdfMEQXBaBkA3OTC/O+BOGq0V58uSzRayJzPfeIFP1QMDr947Anbh7xhvlN+BZ1Smg+McpyYMI5F
nbIc3YB6nc7dwWPKYfEi/RVpDKOtl9XzckyixZ4B2oZFMiVNCK/YjkcE//2xBF/gIZxcLIv4KGWt
J2BicHbXZwZ41F5OpS6AkPA5gMJY2zkReesxYLjuI8xtrDtNWSjddPxIOXKt8R3DuGiTAumLAppH
tZHQw0yVtcYAW/sKi91fSKLZcMdCWw/tYcg+FK2XQEA8mpIhOX0PXKyOILIBcS9Acab5sIw+oIx5
8dvSmQD237KougJT7hYJvJoS0dv22lRlsJ3ZF6gQT+qY5xoP82zO4ex5tAI5wsG80KuWTGZWUmbY
p6Nbx6gE6cyzn55ilLkS2agz3SoFq8WREvHF3dA0Ie03OZ82aR73w0iMGhC9wPBv/tBXb4d6byLq
V3vBhGverRST58NvvV5tHkQCCygFtqW2w3VzHoV6FtoaW4SQrBflGWRrz418UPECB43wvr82oZ6C
P9YFPjVohl+XbLagtlmrruchzSLu8/hJ48VfyPUkXyOdTlJBHp53iQgs5YgVOYzQl43uTo3422mj
zgi0ggcS9K0s8T5ypxqSSwpaGLQmSCG6Szy7Zo8cmd27re4XxhjbAvI7AV1I2/TqhgVIAAGPV0YT
lRrf6M/dClYPZEZzAZV4N3NnrdOcRVWtd8aYbMP3kcOxX6R4zcciXS8PpGzi1U1lrpfI3C/+3xjE
JeHDrx+wXuJUpsMNCIyZeGyQmXrUlx3mA2BFoEMGTzxAbCPsF4nfMmfJ2+ELXYb4byxFipw6Ub76
blGa+7uKiql2xGpywjcXXmEg/JjSguooT2Bs/XLVwxjBj8TGDSw47gJ6FN5nKXD02tKrLoEEATL+
7p+zeK55JGmDWnSE/MuERhOfzVyf0aWQXWMAWTYoDvv93hhKA/OwTa6Hn+qd5l0cfJ4k4rstsi1U
jaEtVwBrHeOuBWHgBu+9da74W7uP3C4WQ3ScMISyZD65vxWWQ9xqIlPABrWDKHB++A630Lj7wdYC
uASLB4zsNUUIdDdTE/YoRq5aBokY18N0JbCFkd0ABp3lC6j3EZbBOkBI7jE6NjrmayPLcABkyXof
M3ypVTd+F28PokfbBGu7/f8NL0lggylqxkZt7COVh08P9JpKHIZxcuTqWbWzsiwxoTzv9pW55gtz
yYbfFzhSkGn94Oar+JmkbbFLOjcrOEBLtIHC242KSChR9h+vTyu3wivNgS9ai7PgyS5Q8BIZpTjX
yUe291zyNIhL7dmVGZDa9Ma7mDVLQp9s8v4zpTowq8bwFM8Dts0wmkEQQes4fq6Kgcby1s50MlGU
S6UW0jLjaufU/X7DFm+4ug0h+lfplLqeVnVfR6ucSwunHIewSTcwcPRu4VQX1cwRhFxyr25meUxt
axC23GOFKmE3lMbqooLoXmMtBInBMvH36rlmqEC7p2bauCeMdnQpb9hA50WAHq+d7bHNVnJXL+C6
5KmjQJL+YMHViDh1DVoL5EfoQ3bhOcoGyjdqfyfwKcbYeuT0STR+0GuSOLwYN7RjYyAAYjuC5XF1
Xhup0oBoRSDUpNbmmv3NhqvRSe4RabR86WfCTKLHu6sMIArU4x7UTHds0DGDEsbgTLTLbokMYZoB
j8PR26sGaUtsjVSH8fT3Mzy41xUqVNxuYSRK8G3u8fPg+cV9kOwKwmxj0fZ5OX7ZVbOeM48VjwAH
qiJzS2/DJBFwk86UGmLMEcsY9OjJuGtKuODI4lifKMzw/tCN/DH0ClZTqYJIihlNJ23w5upjgeRq
yn9gkrWarSUOmdXjejrIg33AZDLwSjmxrTovyoXluhgWshwKIQw9GrI2jGAKshiyrL1HzO9u9+Xr
2XB0Cvx1AUtXcLhogSgYAM7QdzJ/DZk0nIu9PLfdHug/Annyq2AQHqctsLmQZET9+tIlm0eB6k6G
F1Xz2l+FwbyriEcQAEYOwf1BekhWRJCvEPSEd5Y9oQrqeLgRjART73h6Fs3sy6Tvdp7eqLFsyOi3
Wg5V062+ZiAi6Bew3DV8UgpNh5pqaTNmZQRYUBbBmGV8E9Res7bxQH35tijUGJDJaWG7/+ZA2s8x
7ZN1NfooQBkSME/lfZ76xAllZb01AtLWOJ8pL2QbyI7JzLxgnFdRCvKiO3Su6ic5pLEBK9FbzsTK
2svpUwQ4ppjpZ1EhVfrg3288i5JXBXjHbrgI005Qwcbyp8Qdd+iO0Mvc5sxkIsz2+PpJ4QvgUfyc
YDoNOiUE6rKpLYESBHxmi8jmWrvxJg99IgEEn57wE9TRTCpUqCRnlQnbsi+qoKGw5GKCHqOCQu8m
2NLPtCRtSzOJXOpdnpcvS4kiQQUAEN9vohqo/yuCJSZAbesH2LC29izaBtOuB+L2BfxCjmofLazO
6j8YNq1+OhskgRaV5JvGyalWTcEnXcZYfrJzFsZ+eYsD3/GDFFHh4UOqxNyatrgoE4S9egV065NU
hJdPZ/EB3GfglrvmeEdCpuHv7r3h4P+LicPJgsT++kSgGn6KuDG6at0o0WTIAGMCrSr2cAClFjDq
B+v4Aiu+jFJe2ouGmQ5X7lLbsGTi7cBoC4SZVgYLxyULujr+5Fdo7FseHHB4Uvo/I992PwrbIC1j
nZvYirfD0b8EEVK4kseZfMkRTXppVPD8+rKkODqcITRqQAMu7/0IjyB6YSRaoafZlgadI70zGq8N
oXSTSaa/BXdfRBcwAE2wOtt3P9HYNyJPL+y3LdxHMpyy6dE0gQYo2X22u8PR9Zdn8zg45rYLnZc2
euDXl2CrSiUrboRoxvABdytJw420kR5HIu08LIesUX8k1xrzQLzOWeSmGgKlYasuqFM2YoS8iH7B
pcT2swdP+BZXQYlyNhmTVJlAAnYALBQizPACSD/D2Y8a6t/HKYXEmB2rnV5IBEOcrkolT8U0LLZP
4pOPDmcNAAERVRI1Wz2tV967d1mqvgOqhVLoAOhb43NFKkAPFUzBraVid3+FYYt0MbtnMaQ/V75p
IGXCPfu44sT5+6O1Q7hgAp3tjCpOa2sZ+My/GkYZyWFsvSX7cbnestIc7gnz9I1ffQv3MmqPSXdn
nYhZEy44hjHb9oCewVIDfYSePpusih9SbAgwQHpZ5AUBDNfwMI0kExH+lfz2kKx9x8LEI4P/HXvY
raDuOtO5NJ6AMXImErQhOpwQ1lnG6G+UHxwF7jhXyz2SweIm6061vvUmJW+uEV00TDIUKvERJ6Cc
RnIGE3anWAZyyuZwQwemisGvSIc7OscmveVmhl/J7ZwWJaeQ+HcriFftsWZl/LeKrBcMgm4J0/df
8kx5LgRIvql779fQv8XlwbUuJoT7VqWG+/jw94RQrS17Y8XiYlm7C3sDMuHzxx0dN/KDq+SZDa8f
/+8K6uKfZo+DeO9j6gENZiw7NEhVTohU4THLuIFivDsiU37/REJArxYU+gTTPAOpixd75tRjIEq4
fRSeZ0mFV8fzCRx9Ash8D1/6Z/eUfxreh2x2uv2d8BNw8kqso2tOefJbgleQOlEMD6yuV88svLg0
CSH7hKvbuvwi5fjNSz7iUZHl9y4e+BQuvQ3aUz98CAt1blATrRlP8BRVhln+YQnnazL2WzLts45h
Rys+UKBfhrxejHRKr6+b85E+MAjFFFK9r9hHnEcOKIlYE5zwOM99YQT0Laymtd7/ix1Q+RTWvihJ
ESo63j5j8gu12VfkyuYV9h0y2zz/B72kWXNB/1q5Q8dBi6Sgf1HnxI6PuPMApVq9voMhsllxR+ZZ
1T/k0kEeHLtPxKgYIH2M8Sbtbaqdryb/NfKUEnpG3FTAxuW0z5tVj8tB5C0nAO1PBePg5QQmJJQb
Dy5x/IOV8e634333gqQ5Y7IHx/u6v01sHbG0nLbs4epkZiuUWqlQwO3/eirOy2cpcoP6SxzDKNQx
DNwOkF/Qr0wAodcxJW/NbeKXONc8eA3hI5UGprlVsfKCS3z6caJNXqREEnF5F+wPjUvOiv5VNGmE
ACAmGH5T8MBADMGNwpoLK+O8sNVzfRCvbqakOk26A9V7yRGvMdOSs3ny4u+bMzJ+sfMDIgdh8Oue
ADsW7uS4HRaD7l30GmrG46jN1YVBPoNynMR12del5zbScoL9vHC5u4l8Y3cws7PI16AOrjh4IBR0
CKAinFwYLoFuM0c03pu4wAuskK2EUYdNjn5sfWxgbS3oalClO7aD2QmNrG8XBAw/14AdAl5rc7Ww
mTFJDhF+ThWXl3v4nvnXpUJPKwn7pMmqVHEB0UX8NHHnMavltpWKtJ3tkTgV2uu7xtQi/W0UcrwH
RXHk94uilRzdVbAg30kjQL2Xi9Yxq7tq9NLDSVP0oVzI3lM/n8DLRi3aO8649m+YzpfIET6pGrAc
auvA4NGDw39SYZo1SKpnDQ9IKvnOqRv1BpkPF/YX3VNYNSfXx/XrR/UclsjA1kQsIyO2dikKUvj5
UvRWh45NDm9u9eje1/RZ6iTFRvXhVHbTE7jwvSOHBDk4zx6RZS+jPZDlxdT4i7eZjBhtS0sWp4L5
Ut8asOzHniNWbOhdaXJSWBhHM+aaA37Ns6BUXwxESGmnfd1tLgfzSujemwlTYi3lOIlCBDwQADXs
ptdndmykfEU/bao4uMLhN0veAzZArDOW7YaM0rxmBZXZvd5mNxxkgs442AoOQellEuDnQ05Kr5In
KbcBQFywg4K2BGeGz/aWfRdeEeEMhPhWq80m52zEuWmTWp2mJnZjjdwxE002deHGGyuRPt0n+Cxc
Y9fewW7h76lEUPKh4O4NK+nnmfjuIDOgpTxw0ugESJGJi9s69faFivGXZZIDrxhR9RvFj9Hd34OG
wW8pWoAiekdWGLd9mqjx9bHCmRlEJcExHrRXge9JahszSXOwJVpj4CGMQZbDAnigow3AXqN/bq2u
wMuX67hIFWmvSbGqc5V5F1lCYnWHokZtV0ma14fhqCY7CuqnV5knJgW6j8Hwd9Ww0/4AUFR41CRj
bCKYIoDeAwhm3Tjs49+hQPpmKrOdNkqnCwmC6CFWG02v0Vr/M4TzfKr6HuxW+9MSsTVKfUM0eUQn
MzmwIWnTATDjB9yD/aFAbwhX324pcq3SYTZbIqDiDPXWKic6QTuIjnA6BX7viaSVnN2wYUuk90Ma
jd9JEh/F4Oz7wa2b5pplqqC6nOay84d9AxSVj7xOCIAE4+a6T5cIhYkrWVNSdxNZT7oissodQUlR
3On5kA4lQvzeWowRBrVrMMsyFogKi6b8BHbkSk6YUOMgthRQFRVeVWLPeboIMHc8idrvh2SxFTMQ
KWfkMtR5Bsq1GlJAP+oOtlro9xvgpc9u6ZjTwnEC4yC8RiquPKr/uw/AEwJHJu9ZvweTR/As4ZaB
uqltPEqDCpaGuT7V4Kc5hCLBc/59BmywD/Hqe76BSdFy8Pu1hPcnYCgKTkP3GHF6C2NiDM2G0HI0
d1/1Q6Hfgn8FqI86mRZUT2lyzMdSCeelWKH7MPAcYMG39g2QOu/YPQPU2C1JMJCqeYGjhRYguNSS
JA8+255IynjbE44xPEoSWnvZFkp291XdmPMDIvrR5x46z3255Da2QpNU0lgE2NCHE4JBdodz9kbm
Y+7koOq7ktVpy1khqhA4EYqnvA7f/1BNd6aBYRhuR0In1R389M+Oz+s0B30qoBomTGJzPOyCZJay
oB35dHgxeAi/7Lg8ugNafcCPxK1RqxCYTHDXKcc/cMHhvVfTcKRo7E4wYnCXstUhxDtc3tSZBlsc
skhVhZkbmlRvGFuro40BdRCS/hGCvhaAIT44JgS4j+lbjUyr6jK9aJPND42osJgLMcuoFZz6WNUd
NCbIAYxnWbEj+iY4JVDbXNvx1j5wt3mOTQBgj0/y/dlE650ehJIgVHuchT17VlctGG4pe29AK5t9
sj0xekGOdFvd7MXn5f0LyIqhAFTUpLyMrmKYbEzuiSiNMcAsMkfDEGvsErEFAlv22r2VTYSPRZfa
20JJWciOAomLdVXK8wFQNCYJ0DQy/FX6VKl+bX8UcxfLOOIeiTN+GFd7oChyR5ARO04QnOr/wFVl
kJxOLogRp51kcPrGyT6PDsmDL7ADMKt0I7Vn7Zf7VVccPb8HEZkSIZVxVbctsksVKWxEBTWhwalN
diqfQ8z1hRrULwZuEGyb4Hed2Wtq+i+wbu3ROA8YIQkFMSCcL+oRCYea/eb72j5U1qbWZeUY05Ho
6E1vajEA8hrTfTOmeRY1e7w7ws9hcLLd09zdr73zgvdnsh9Z99qP+5O6BCeJQpl6K19QMvGJu3Hq
SuZJ4Mo4TXlnqpBEALMgrc2Ji7l08SyyNvW2Bmb/3myO4lKGKKs+F9Sehi4FqkN8OxTkBPEKoIK9
U15dzh9pwWzLPkydZ/g3jgaBw5Susen4zwWTHbNXo7tFvg0kmF1mTPu5Zcr9yQos1NlsFyWQgOx3
pn0fLxMYBWvCmEoGweVNGWP/ud/pMO5us5OiL5+LM6if5Uu2dRCxBiNkClgL2uAqhox+XZd7DQF+
iFYEOjdr2wfaxGsz+BmM24TMDLv+jwN3urbsds3dwtzWb6tKK2riygwX+Y4KJ9ozB4E9W6VxMZ67
YhL43/wJOw+Ik4MCrOgrXc+B9hC3tlU8pPyJahHngQ1iw5il5AaY+1cld2UzMf6AwzwEaE5BCnxk
s2tKV/NtVBOK4nhuO6sckyA8NTRAaE7E+qeS07Qdnu6Id0cft2m9gbtUJ59ykV2sYZL87epL1EgG
8vM01gb939Us/tJTEK4lGVoOEAhQlrw6EYFGE5Smr6ZgbB3AAAKlo4Nk/esu4V7q7EY5EdIdn2Zo
goF7idoyw4zvYa6q24yGn9JkcxI8Rgfota6nfgG3Ed5+6wLmWppVtUJHOvvYYVY4fkG37PHu6UYk
5HSfRFaYgbsLyUki/q+FF6qKkWiagv2S7tlaGy6u5tyd1EEZIR2DUo4GQZKEz/Q9OhvgX2xewv4Z
0hXdky6iNj1pZrW0CObX17fms3BHEgTlCNIvhbY49J4q5bxOY5w9qXuUz8J+/i8wIae5Ex+AA4BX
P5W0FVrM63xlawfXYq0HpggfKuVJuVPkeP8fFKabAeMKs6f5glL9P92xd5Naw8yk6FdkowoWIV1t
xjhAy5itsbItxUnHagpbJuvO0TlKhEPZ/vIn304SqS0hJVUlGD+2HHXDOGGZKrk7A95vrKzHYOM5
DBUNKd6MjSiUVAjQvlbEr66N229/VbOdK0G9YKriXofU/RLoQOgX5gQ5HCgUfZd/e550coSOM1r/
hVaR0HNy3YqwGu6RfJ39pIIgbNum408AqdaervbgZqYzXO6vp6a813cNOQiOjYwYxCyPzXeeb2Oa
0QDdMALgUX7mVjssVmZwArFEpN191osmTXBC7mhk6zjOZUQAzdSEo94iHK6pE5tYCUN3Q439sljy
hUOrNjENFP/uyrp2Ki3/c9ndKcPVYhGeUbca6JxRSrlSUqBHpspjmLpw+e5Q5nxk+NKT8BWWNKQq
f5FJHGeh1f/HuMDbeEUJGe2Z5Bc4K2KxhhP8sYIPkQ/YAG2C3Y1fHmev0hc+vdo0f7lijMcgjpZ8
xgiup6yXdztjlEhOaXcrX+CKISk6bFaPE5fXcgjtVj0FyGpjaHac+2bx0o9hQiHw2cJpwi25Ngux
bTLx62zf+59KVQ17mav7tbfaRj6vZ6qm6rWt1AkR19ThJPJEREUc88jQ6xr1Dxe75rdqDcXZdc7h
PJdVXyyRu7Nw56EiCAYxzIQeGBlVtTkSuGJDZaO6ULOrOf2TwyMfjwzY1mxDSzfm2nAYR3ovTeZu
xV9rN+h+KBfbXlIJH7R0Dz8I0kk6wKBZTlSeSMVnLG5eqrwBb+Hqc4cERjL1Lr2H6Dj1whgNwDTy
EPaOJXCCvsMeBMKbLkGG0HVigzeyxVWPclbQoZW9UHsEmpNdKgjzj96PJQPABkaWsbRHVMlNAPRF
YwI4fjaFHJAWmf2semtDq8vxoB1yHj2M96A5tKSIj701y/KxshhMNK2CC0E+sGPvSOdJOckzVaTa
mVjd1L3jzGDkl7WJT3LMgJjAcxMOt2Z/NhIRXgrixhTT/gPC/Zi0NDmtbxyz7rAg07s2jtox06DD
wbDwUm6o+vWflUDbH+KC76YVyGB4RQ5PC1xiwjnraO/LHR9rxLJX3zx5/DKd5vP2TEudcBsYaofd
UVa5RyA3V9gif/jvYGdrS9HGakZRlK1fZsCoTtCJNzYF9q1d5gZysZjdw0N/SAnzNTxaBcxgLHfU
qU/gRQqvs+knSz+p8K1WLw3tOd7cCIiIxuPYcybv4iLoa1Ribvb7cUI4Tn3VK3Hs2oXDTPBCuQvQ
o6xc83doND3RI3NCFoZqQShsG3NNNnvoD7zEIKleE1T4FTlLFc4X/B0S82w+fHF5m/X/Odyr2rP7
061w1qpJLi26g+sZ756BJQFxlbvYNmqOeOfsdkQ9HdXLwrH0KWw6OAJd7euq8LQo8nN/9HHOy5QB
1kNvoG1Hpv6FvPdksBTQ6pBtj1YNRfPa5uQM2oSrHNRao/C8mh5XEhQ7E/AeHSxYG23FVsFb+S7q
3XKZmKdp3YQJziWUEHiQbmxDoLw0hqKGa8d0S9WpLYnMd8CWjMn/iWNU7ZhpDrq7g8uV1eRQ4QzX
CDc1wmSGKrSCbFnG8XDQSkNtMO19DnXXmnqeP+5Qo1FlhcUtXuK7++BCj3DyDlCW4YunVXM2AYod
gcrB22uF+OpJPhoH6oheB5ZM3+/ym7eRpSUiUcCWuyfyIt44+6iVzXvORYZp2uZw44LOQKh9BmJT
YN91bVa9HIDY36xdv//pluYuFN5t3lA2cXgPDehbydMBIbfUhARyjB6J/G5mr5DmgVxjk83bEyEW
qs9HvTIlylUdNQbmLJiaf9DuiwGyu7nmX7nN1NdJ7ApkjFzkcL3Ob6HvhFPm7ybT++BZyW/4GIAQ
Mx6eLGC0RPoyrCNz8/uI8lcVoeTmufIVRZsS6pGnITqtrgtYEI9YnV4JRiPi5erW8jwjN35do8Lf
0fVRz5rlBtVIfM2W/zj1bTH8sjojZncSJa/O2D6Mg6RW2nnIr0pWFdwvWHZsEoo0OuAy00IKzefM
n3l9E75W+Awor0dn8Yr2NRD8ZFX6TDELh4DYjcwMlNEcPaoH/rYUfOXZp6n00+PpI7qFG6OlGpjB
cQoOV26Stcc14YVGJJUtjIQjUC5XblKAPaZADRCi0uthtiLNdjhEWIAxwmTRDuOBZR1pxIJzue8D
ngVSRSPGSgDwwhBbaStgGkVFkOt0naHea+MRhOcIrk6LHZeVsc3Brs1OX8dx8AlHCv0pZgI/+8bi
BP+RREuN+IdyJZlxUeGe/JzYgfmG5cgu+ZBD+e2D5tTjnvFxuzwoeybdKF0hjyFAGwuAoam+XvXV
9LHsXRFWkCd982sHRZFA8eO8cjU9myruKc2dCrVXeKCVAavQ+JljF/E/h05o7M8l8ELNduwFehl4
0NkJ0Q4POUMlO9LatQpcFZUKM+zM1zIamyWwKiHut7DuCZVJgFYqFLjrv5FbWkGcocCq/CH/d7XS
WVWnExsPQvUDg6+SYrf8GyXMvXQmO7OyVeeTUtukWEwhbPeKfPdrS00N0LjfCf85/xWfzN36+S1F
Brm6YAWc/bnTdyPisl4s+HLkWy2qN3L8tBkUncdKrt9pHmt5PeVtoHwWA92wq2+YV1EczKaY/0Na
xuVMdPIyItB9V/z7J2cmURYob6p3ViyfO2P4aGIKvi/PwxeLUKK5AN4WlTTucSE4JLRaxbpSUAOR
Nt0FPFivBcgDVd4QyIKB+p5uv0Q8LEHJTJDwzaboTrPWlOQgGIYePoalQBDAVa8Epn1HdJ8J69y5
nV7f9d1jez1M3+nmbM4RtGZqJw5OHu88gmsLjRSdDnVWZSMlo3vK0bxORQgaISqnQqtyFXvkqSD8
eo45N5uV76McHM2Soj3HOcvkOxzOXmpuT8lnhuzyHiAK6WLhDg3DTGaMMtzAClDpIHk6SkvE0fcb
ykfyTO/F3Jtac72OFvAJEZLj0hXZBM7x5prjO1XqVlW8sIwEyyPl2s16PK4+2VELaY9Oile+trpe
e2mYJeJpIq4Y6ucQQatws4LoR6fSzriK/5qca0SN9t4mgacFN/ZVEO4/KVfr+LX/Mm/KA41h9Z62
naS4aCjI3kmo+cQSuHzGxM1mp06kJcGGD+wpKOHp2gctPoFSmbYOBVCGFpodZwS5c+rnMpCEfs5r
f+K/rPV/laQB7McQ4m7lF0tsfiBQuaMZn1sspHcPfDFUgh3T1BNr9d7PLSSt4QABgqIU1M8/TMwT
5CFAZR0RQNTlrOtMiZbPRRRNnUn+RwtZ7yGQJkAQuIL20CJ080Sb0WVn/xpCvcmc5wcJwPin1QNU
YTsZg0dD+h/X5f7E91mODWCrmOrZJo8UgwYk9qWgEljsKNsLov+CHIsreUiZs1McoXfvSYdmlS4J
dNcHMgJo2zePc5sRTwm1ExLtqPfYQVLU81I1HGAAcwQxFxEBXXNXd9/hg8JS1ilJQovGAX7cHDZm
iaeiCph1cSO//TewGn2kWN7MRb2tkyGvSyL73IE1igH7iUnGw3lnkqpSW9ayNdfho6YlPSmYj+yX
IH25CSFpRelVgDZSNfpGXQz9mnacXQxqGEiS1bI9/o7+AmGaZMc0yJOZroVnQhK0jfSiXRBl39N4
pxZTDaRgxmONo4s9TxXwpGPENPGbQ8WqK2g3ME5e3pb0zGkwlRuj9itWpbWhOsxIK1FhvNUmPiJX
kq1b0wsjC+Sa47Ur5KtWSf53qjm0/PFLprz0oV4JCZ6g/T4ijcXTgd9taQpeCsq56Hbl2wfh/BTs
qMy3Ut2KFzCDR5CrKCixGDljTwiYyGA/qhw9sxC5b3ZucxXxDiyiSu2ofcHKLqcJuIZDhkGN97sO
O5Ti/b5bfC4PftF1H01rGyDQfFdimBhM21sH36LzDR1t2WbHhWIhcyVYgZvdZbUEQj3m/l91wbIY
4dM+2zh8qZPdGbGlCnC2gwxmFwAyi0eXIqMftkh2YW5QmGIxIKsJ5E7FVxqwHj2Wqg+/mZyiaOxC
rZ+0KNd6M0c8ixkDh4MPO0/FUGqowQUYrMGSE+J8Hqw9f3Z73KfenLOxWSJk84Qz9an2AciF3H7Y
fHFaLGdm/fy8x8H4ckU3gnjQQ0eAf1UWp7+0He8uP8cJQdh424VOjoMuzA21vsAtaBJpUwAvbGbl
OJoUJYAxX7XYHDWLxIQtMBhCJ5NRt4gf3CxuLJGd6rrKKsD6NixFSVF+5i4ZSFZDBisNouuf1ll3
mX7G68h9MtRM5M6RT29FRMx3gfhmNvHTL1u9WehChJ1WW6WwjliqJ3tTnjZOTRVv1r0j2kDp3PNF
gYUghlPM6XdWLU2q/yN3ZKeKvRMeXlWO45sqD34O6ArCTPvh6Ri+ByKwme5PyXk7IRJeEK2JzdWa
Vm8K7+xZN9oDB9+gAAiZrau35LQFkn7RyZ5DsFne2Phq8ovhKJreryz19I1qDK0Obx/W+fQDPRcq
TIzlHeNt25ApVm8TlYzN5lX+UORF+NjOq5CRZW00JoYFqeMRtaZMgg4O93I0qFBMNstpsSlIBgmA
HIQF8I+pwVxJCLUNUg3sLt4JqbgWANLpcjdNWEY5ck27OxtP65Zb4T+W43nBZiJJ6bPHHjIWWNCh
7uDFKJnuZvBPPWrPUiy0MdFqqCSBh7VRysBm36qfFFk7+/li8GHwvopq/MalixgCqeDpsb0HHchy
hdiXNLhSpyZnNKl0eaY0r1F6DeTR6UYDy8flLymllBW1hrpXcx7zMHXbcuNNvJo1Wn9CiQKXHzRA
a+6VzHa1BHgeNA7nH7+tUHLGiCi0mYXHccwe3nm2ptlXQwP/dbkhr5cg28jpCfJ3tOJaows/kYkj
/I/WdTwtF/beE4xqoyTl+ZSJT2H7ijKTypqybLVB0z33nKxi/hfeV997WW49N9zgVjf5OJJplkqa
WmqWXOAxhvFM2laJDPv5jFbVQDQYGMNdxV3Z4+lbnlrwLFrCxiKiHjmHgQzGWxxsIZsJ2OVUkCDK
cYWDTtwuAExKUZDwEK/2mOLklD9XzXjRaiQPL3V8K1pUSqwQ1ptAfPluOHybQqzTLXKwfSgPfPMY
Opk9JCiINwat8uja2nrkIwEe4FlU4966ypBxlFL1gS3+HwCPFnGpG7nxIuJIF8l0ngslYSP4NJZT
p2b9OUVdusY+9GjszDJK6ov4bvLIeIx+2ESibnW9/HSKcHkEyz/whiryw0WJbR14wPFw4jNThiXS
bNa4Y1qMpVyH1u7US+xIHTIQJJoZWZkT6y+6bqxFzjtT2FYbKoyXfhweeNrWieykt/qPOLSaW1uB
TGytvHxDGXwa+3+iR/uDWYM5A7eY1uKS5i6dXI4GJ8Jn8+BTs1UH3GJrwTIYwj6t3FtfrPrKRvem
wUKIG1uDN5Wr5R5kJwUTnGwgK7xDnrhzahDG8TbdVziNB+6NjRxHJeNGGfiLciPdu1ydRRSIODk8
uHYhpEuSQe+iu/FlLlC3toPHPypwunaW54twYYNyticvkEIwSUmrCDsN7EQEYTguqMqAuAi9Nxaj
NYwSBKcEPpsqQv1NbXT0c0g9lgK9FKajGnA53MMvcPuIdkLK28wJLXjkkW6AXr7LG0l+aZNo+4t+
smcy77z0+xeKniJT0ZlnHhwK0bmfBBpn+PtonWvhwDUIaepPAKwRKZhDZMy7djyq80JZ3I/phY3t
7tgsGF/ZxKgM06V4VYsIVBhnWiG5aNTJNd0drvgMul3L2no40Yi3Ct5JPAutKLAR+EJNBYVUb092
s0XVuU3O1iN54Z5jU/DDHpHLYY/9HoBzj462/se/Wy8k2CfhR++CfeUU7vYtU3XpKoNDS6OwBaJA
B9+RXMS52jyYBd18NvShmi1e2rIXQjiBCdT6Ql0PAMe9XQOr9UsFjD3nYfYLemaoXfnU4mvmEprf
uIWEp+HP1jKtsQRl2CgLZyod082KDm2W4cdxjvjm3bHtd4WlqSkrEzTx97+lIHyfDowBFGgkStZN
liyyD7Y/73R/8Dm4JRGK6QxuvfVJ3sK/oxwPCBOdq/mBPohN47LuabiEAFwEFTrj0ECk76PxGE8h
8ah9KNosqIzZM9O39hyyrratI+5VTy9q9BfnhqV6QxaAtwSIr1x9QAHzWOx7PoV1hmaS4owJEkbD
SUOUY3hkofQNWvuE+Lrm2TOPlrQdzH1QRK3YZpeboKb50pVjzVQK4VnBvy5oR3ZUXSwL+VnWPepV
5qt8bHLt84/RRfqz627UXxl7RmTbbb66kCkQ05b4V6tRIacrAlbm7BbmDhx/OtkHm9xgG47yfglf
L0euwECFHpUN8KJTlD/2olRRodhBDr+yrwfUG3mZfNqnPIrZ2RV6n7X1Ts5Z0qeGOZgSNA/SqiMA
c+sCvTuSA3hEhyxrRIwmqZWwHhZdDR1q2AYkcwkQcGihFvnHQh84K/5SQsRTVnUnY0bqahe3hZXy
v3CHjKqZPvGKOc2seRjUBYIYstccAMmn4JID1Qz7EqBENvXYJ46xQR16fB7DvsMX49VUmBWqXGol
5kNDRkNNTb7VIWc7M0LxvjDT3SryWiX2xYJGU31VtL/dqXnNtJo6iVgopOoWVhtUhjwB3karvWtp
MkPVXIq0xLS8bo1PkpQliH8DXN3HNK0Li+xp5Xms/gUbAyZ5OJ9kuukPjzulltq5Xo0aZrB3reAJ
2I80foK1qhV4Ubjm2WgXuT28llwuUoLVzL8JWShBsLyXEler9hUdUP3Hp1MHWqxM/nvumVfWJQu7
v1cKsKkebBhJGKi1HMwAZoHBVSGXq8bo9T6+R3iT9gx0gktr7SHD1gEoevfEel4Rp67rgrqTKl4v
LydoRGYr7Itc4OZrDMW796UlaBh9v1ew6XIndIFSR/E0YhBt6k1mUt6YQcqneRTDgZoy5LVf031c
Zy9y1KJeLYuX/qIHGSFT6sKxxYEsK3ox0m1ec6mB5JgjtBhKA2GvegCEyIMrsuY9dNSyVZYrNGOs
3DKCjQ5xGsZmCpN6YS/puY6bz7rABvy5WS19qiKbz4M7g3aDW2PDOZaHjbhvcJcUqrS4SONvFcLi
ukXsZVz40PX6G81W4nAVby1V35J4eqA6m/VLLOsQtZCL+dBM8m2F17ccQ0ysiOtSXCmL2R+31rvA
TnbkD+qk3pF6Njr5PkuoGVFgDsM85s+LldLx9cI4EApZQcR2Bi3fEoZEn/EGSuxHmkRpuRiVdmU/
fQXlbBM54mYz4Tt1I6yEBRSTKVJ/gnwUPS7qfgPD4NFaARpOp9ME+XMIjlobUCuMsJotUKd/X/uo
KeEuZ0MbXAAQ0n6iJzuYsJWV3j0vvenDKwusJNiZjDC/J7RcfMGyHx7r2vLrZkdNLtN5d8rfL1uw
4yec3wJtoxhF0oAcztpqFvsfG8dVj3z9JHizEiMH9aMBSYq+46w8wXKMcOppaEhIYLGtIviD9pSR
tRbwjru4V1BgAPkjKBaJ9Nh7cywT5+MCgrBVnRpbGIF2G9dq6mw2SS+k8vs0D55/FZwvpRMspWH4
S0uMT9eKspV67efR4zYXiwUin5QVw1JyN/MT26r/tE3VQjD2csAGkNu9kyqfQyYqJ+3uzemBudJm
jNNjg3elo7s+YJZFqFCrjERJ5UPsdH1vv68kM2ueCvOvoxTDqZqsSlaUaqOo2+Ac64WLifvbw/To
QJHVdl28y8pxav8SFIkj5geHUY4UfeeydGrWaufdw3mDSDI5aAaUtL5XiD0QhHAu+XF+TxLIZgbT
82Wx92xZnAh65j+C1qjSMCXWmb/87eXO4/SmW+5K/FajnbwLqTnewsO+pRt9iPT+hIUrdFoMu3YB
caBbj+8P4YGtsE2TXZE9lGFlCxwTnTEIgHRPcuibrHinTikSbJrhz4PiBdowMFQOtcxiFu7lOH/8
3wVLAoKCsQ0K2OzoIhsTXRlXrA2B/+t09PKOEHBMOC9/uUA16joSn7lUA130KXAWlrZTlemWvM4Y
h6tBr7c4qW9fd4QJWGcI7GdE1OVGr/N+lzlwNnrvFp2Blxo4fLHunYJLduB3+eIxfCSPkLIo9jem
5RbgvnULZ7ytI/Fr0H9Hh/AFA21rz8NSTY7HM8kiDY/aJEVgdzx9261bASRTfhIssT+nAfD2OdfA
rmACyBR+Svsn3c5GWq3uFnRLNTEAwnBn54z+2ZDGfEr7Vjv9qfnnpQU9Oq7iSgLQL2FId7r+Fe1C
l73BiK1P9Tgt2XeFAuQL8hz5ducX400vXqAGuwrqWuAbuQNipsrnBb4gcANxd7j5NhsOhBhgLkEY
ikDaFg2p0KQyo5cNL8KOfD9kkeUCd9eGVH/deL04RauAT5OiSgKdYg2i4wtUslVHuCSo9fHQu25n
XeOXwpzRXWLManPeSNf1ilg3Sh3Bov1rRanKNKqk5SyUY6Fl/aIIFOpCKzK/JkfP45XMv0hrM5x2
xZ+vCcdS7pT3jXSkj49M4OkVFSLwWcQvYLiB49Jj4Xjo/Fw1o2qujPbdZQ8senRy0ytJwg2NuAcH
hOmWL0zJSD6SPxds0k6KPeSret5xMUGSSPUBy+o9lYEvu7X1H6k+qk46POPnvVpaPs5cbZsytl48
f3SHP9Lt4hftoUU24+/+ZNkYOgRp7iz2mXSPjcB7p4fhS4kNy6MuwfJPKOQWnktRRXWi28TDnk8C
EkvOsuKgW4LM62qyXiWRdzsScPLmPcMtJmoze4xBwgstuoYvcSU4MPvaVn3807rL3Z4Nty+e58Ay
0mAORJNEDuTq3K60Q0M2gHpyfbv2CHJFvzVMCxnzUtLHGusm8HnC2qo7gez3i10bn46sbJygtgZE
ZgUi9mXxq1j0fU2e5I4j9nk9VwJcgOH/OYOwNZOxY+UwwQrfw7LaoBHq7pGmY72XRmMbbLcr+49O
AZReW3f0rq8AK3gNoMUV5O7HEYYMwzGe4MlysJXEi5ndmLi8M9o0udNKc8+yz69NN56GkQA1G7PD
ISRkcHIJDCxvG+sjweyrcm+OB+FxiAyBwFZdvVKW7L2HOtJoccrFAipBG6hBHVuV9MZ4ICN8REfe
Gi9GTLOkD3SLM1um3c33132ZlTQrtmMpnwMD/V1gV8ftqtRMDO6pal626O2mjWMso9BRrHBp0isR
xgG/WCUNIv0spSWy/HlqH1E2s2KZuvFcbVxajzKomA+2Oz5B+NrmaFWoaVJYSbhHqMrtIenS0BJM
xeSxjuODKKBztIoz4DRUsclSaNpy+HoOh5Ptwu247Oj2dR1FtK2PrKsVGFD1jQ9+D/GWnT/V6cZz
CrwtrVMwNpsL1ZRdr61BIKYIAt6ZQ2xhu7NPJiUpOMhnYpnwtZFMhhQHKLbkee2ueAWJHh/N7UIy
kE2MAe/qvafqhEM1CXU/bvzB0LsXDvy8ShPZ5QxxBVZuz9CXpwAYLMhaykMsos6pBETsME0KeoTJ
1UlJ2eIeew3RAd15prIB9vllamkqpDou6cbknKAqPeOeXj9H3yYPol8FPX15Vki5Sfg6o+JHaYoA
waWklROsXUClsMgrWS70AHYe1icWE+YVl2EMWwiShhxDgW6YA3fdddHulu0mj+8VZMp1ExbbyjA+
fXZ6MtaBxoQMFNTgiCKKsouycF1I3uhdFRaevMkFPpNW9U7ombKnW1Yv6Z4nzK8esjC8b5hdsUjK
FkkgKc1BRHFCxRN+kPcog21+q/SwbyZUB1yNxGj1bDS3gA+JuiOL12a19pnSOZ238rOis3N1fQIs
ljZiC+zmgb5mRiBbBKM9vFgZKOc2UCjsrNzQ+QEuYYyZ2kUfvyduzhSPkwzhpES0KhY2ZIlzCNi3
b2EOcAoc2TMpdqHg260cFra8n2X/373xCW5hHJ1qVi9ru8YBZM0vc6S2eppvktTZOVZdkjh2KfJ5
ttac+uaj4A+pcMkiMkTijkybJA9EKCQh/rdmAgyZSD3PQHOV5OG7F0ISPGTOBdmc2CShyjlFDvQ0
44asrdFz9jUFMQCx6vbiDRSbR/eoOTlBSmBhyX5THlqwe+osj+fklxwd5bVyMxBNZbWWd2/uxYOg
snsBEucPQufRRLnohH7sRZQL7iy8KzVrPCk2PA5fFumXL4sM7PtQJE6fm2nPLjWVHo7u56WXQ4zP
/aPbNM/XswZJ8xsCR6Omn8qThFDxZAQcvgbMPg1dH+eINNSjUPK182gMkNKks3Pny2XOZj/WrnIh
tsKLAgWh+BLVDFB71Z6pl6wscY0+GlIceKsSBVIkjKO4bVLDYabE2l1tQHkwqOZPIGVGb5yGacRQ
Iu5GCF5ZaElxbAfqPmnDPRTWJqHCThZx5ZhHpPUhcSIL/XhEzg+YREVy+jG2lOFQkbbMsxwF9yYg
008JVGu/vmPWRGwGBYwmnIum7IXZoYSIxk3Y4//bLSppzJ+D0a3G8AIGpQXqqB7UyE5lI+rf6qTE
yHgzetWus4Fiv+x0scCk3XvlEZoxP/I54AGD9WuIVPup8Uevy7mfZDBbb8vyzD8X3n+Olg9aMnER
ZNDV1rdByFJ7wlcmPoOx+c8XAVFoBk3SbV6Tfk5O40rHMckRv0o8CPFc4BYN9BGhJdYEx3FS21B0
MXU3rmKY5tcvR6UEQlE39cPo2jeTW7IIKhQ1TN3HkRydy3LXsI3qPwQrZLSACiJpJRquQBtYpgVR
44PbyYKkhDtJlI2ZcUyH6BU25Vw0OEQDdjTowu9bZ29X1n2tDIaDs6XmsaBFCN36pYGcxwoOoF4v
i+g2dMJbqe8f304Ujd4aqD0Df7UnzNqaa/HhopBId5ne5A/E5oAD1zYoin23GJei1y3h8GzvMbTL
v/T3lXSuUjTPH4BWtIdeY3xtmbp5p3Drn4KIrBysevym7bsbetHwxjbcl8JUp0awKMjHF0xMDKnk
6oUyN/T/t15KaWqe6eGRhL8YHNRnY7Z1bTBaYjT6vJjKwoJ+wD9uv0UabPZtgDjbI+p2tmeIdU51
6GGXZjZnc4k5z8dDRGlxaMsjC7upS37jaiHckuKcWJ4hC0we0+lw6grOy5qr12Y1bE3en4wvSpcf
iqN5wohxTm4BQ+oiEgyG30CTqu5svAfKJb+bdY/TQ1QlZvpk/I748DCT7zDzy+T6LwHgBdWWkQdX
h+6V1hFD9scVjFlJl1ae2QvMYpY923j0t8qbAQ7mi2AgGzmyrVnrIugIsOV0LBkIP1P/o2B8rS83
9Z0Os1GDVGU8QJ6rs7rBvIJEaQLpMu3M+3Xt4VWDqg+9s2QgatoFHgQTiZRGZzGQ3PyQ3kj2j+xD
yMpesP9hXbTZvcGHg0rIOup3KxJuFjsyvnxma0isqvnlaRtUGmmxx+nOWSq41SNtWopjywgcaFSz
bVr434Vex75rZTmTpk5uh/9I1LrDXq0n6bn5AsXO14ydjnm1sdGrCrxGsA81Jd1M9/Bnua7WhBI1
dTyYH3OrfeONGLkFNphzpkDhpAnjoV86KONn+1dDMPtbM+Ez4sgfohpdpolTgVJmgXrkNpaWRk2L
nqLyX+CllVi4cFJH1/5ynZJcFjw6iraMg5bI0TPnLlRilhD/nmDKDCgib4npq+tExa3ROjSW/JUX
x34p5984W1zfHQWC2maILUkhIT4eSZ9gPMnxHMaAPBv0H5WIyS/YSl6nxPw0pqyjxCs35RKZ4Zzv
HRVGlxzHPIYkq2PT22PxNT2VBDM2aRVQyFyojXTJlLMfngDDSqsCTxwooRE9uHAL5lcKjIcxH5YZ
/i6+V5RX2G5J9T7wRSsWOtcqrdwlGGnGGiwSV+OWb6XFPpVRARWtwgJs+fL8P6JdYvX5w9RJcn3t
El4a5UZs40IMaouS5ASyE+X6jKpHuFyEBdEE8OI51m6gxP2oXneFjBXUuslrtF6PjbM6uTQQIKGO
fPUxrF8DBK+vcPDYG7Bu+ZvDdu6Hm9R2NzTmiwJ2/PL1sTYvMp0iW1Qja+rMb/W6BhDR1A2g+O/2
k50JsFDZfDf/gonSAJUZjAZ7lSKFRaiDw0GHQmD98cWE+PrlnPRuzRdEhre/tKI8cByJBt930o5w
PsGcrfXgNd2wUdBmo/11OE9HkLanmHo3fHBsYjti1x44LoSgghCBcXpII1k2K0fKlEREen0kZdGj
HU1cVNlXnO7vXMWyltQBQwkYz5tBO+KV2VQ8XYWOAgLIM1faizZksZrtWTBUaIke2LWcnUPCesP+
F33HXpNrjvYKxZ4XpcUU9fDpgsFA+gxKr0pAjZ/x8KBM+RbescPs3VQqRgZhVKOyFN08CiNjSmX1
jrNlUmvD/heibu4dHln7AKvnb7achkH55D3OT0jgfWj4Ps/T18Nf1a92bY317PxkDZy30JOto3pI
uSvsu8aS+UDeF/iGyLH1cBVnhx4hA1+r8mG9Sb6PZQpRfLIOXUGclQ7Ro5HL2tU64D0fXy21nX5L
ZE2SAtmrHiihJR+ihDBd/3gx5E/tJA8qLjQCxdq4GHpw0EWqtpS+K1XbMYl+t9izoiulCKg9qPgY
mT1OFdBRy3ChID77mINzJn7rG2AM2FxAV+m/SlKJaC7CTXtvFEyIq16hNLlJxhzojLOCPdQBCLLu
qTTb93MytfUo8v8uAojiTNkUPACdUGGA/HMVDf51v0s31XizKhEynzyTPLGVKrbI7+GvckPzkr3q
DvXg8950IfWsxn2JIs8W1biRlKNEFYAXhB/jGsZwf+0W9zKT1ujftzijkfosSxzfUf83t/Dol7Rk
MceG4DiQBP7HxqW4sALV3z99v+nX3NriLHLnfTmpxe97orJwnKcpLfX+6FkcvAoJCyhcW/H1eFeC
wP+ia7CkbNSCIRXCIdWDMAWs6jqvDKaEi6GPme8Y1ZuEDZK4gGXsIlTzWTUx9d4nnyG/3lkYdPY0
HMUdbpB6ejehkA260ti30XVqw3hO8KvC/G6Grt0IrT70xcCPX8bqn6alaH+pDXlyuV//7nqnTtq1
ZbFwz3qj18vvfMaUnQGNB9wkqy5xLiBbdXK/nEzNgujXWS8XotUXC/q+v3qrWjJI2/uPDldMNyP1
wt/vyNP8sU1Cs6Cm/q1PDju/TYQWmzaglHN69YQwiCkpoj+undyVdHPIXpd2LUykHj/LuWZcOK/A
B2zCmaS6qT/rK+7wbdaClTSHtJGtiPK2EPWPl0AeFhg3ElDg48TmalP2SLUtuC8t2S+W9OYNjI2J
uNfjSt+5ceX37PG4xp60c079tY8nSMMf7xWLmJDYHtKUi/tRXPLA9NaG+6MxPpZzbgYic97r7c4l
pjDjBivSUCbg89m44UQcXcabegmkR1SQoyVxusKa8zfLvEAWXtnrsqmYEyuCCtWgB1qgf/6Ysc3O
V512RXeQ8UdRYYEZPhBw2gO+atCwXKa9hChSJxeNEcSgIR2xrZUE08uHII/IR2Fv5cdffqveRoge
6CnVGvTG6csmQKVrEZwF6JImFXbJPkuty2oW6n7azMm4cDR9Bo91uNF5lZ+WIp8EkgF5EdeDxRvy
UWeLH4eywRZObH2dWNxr23WtCXhbI0Ahscp+spXXiZBoJVm5ezKGpevXsu4+mzGE91jXQp2xJd3C
FsWuGOV86DvUxzE1Llv3tC3hN4HCb+u9vXuCTGOmPVwexNlzLviTJ31IvJ97CkVvsx8E4V+i2Cx/
sfQsOft+fZcYzvl0epWfCQ6+n48ziNbKXn2F/n2020H2KKDBUsvjI0W4x/T0QqX1AyptyRThmlG6
B9MLWzyWIHabiHPrxxCBuIheKgdZPD4mJOE7j+/kmuH4e1BgIE1Y1hcVeO1zu4S+ju6Gm7DO7rSy
3WMphRSiep8OjU5/YodOlVqmM35Dl+MlRq9t5iLp96Hxbc0RvTSiaM3sV75Vkaw9eJrznrhQ+G19
OBGLmJFm/gBlKwER3poX4ywFpvCAydNCxIn2PREOSX8FNHebciDDZXM6I4NhHQX45kBjxq/9iJjX
5hAzVI5M8GBV86I40Kw381ZhjrRMsOSaLc81a8r9rKrqy+3ZVB5K8/fsNGK/7QaDShTQJPaq3gK7
DAFgg79qrYBhSVOQ10uySIYZY2tFfdUu2kTG+641IKf+xFBheCzabvkY9y/oijOrFhTUIGk8UXdt
e3fKL6+ZPDx274pcY8Nsdb1vBYmSDpyWOzvOEiLa9xThTAhNNoHO39qIYMS43Rgj7LK73DRABggw
PZwA8Q9I7rtIWUNeENbOni/O9JlXFmDkf/zNECgXTnOJnbvAqHGFtS2os1ts3hhfrlL479FebxuW
CaRjLBSA8JgxmbfL1XMd/pcANcZTYRgs9nxFUopteYTKnKUBic/erDzyJ3+rNPAvTo7a2cnkHpxi
I0MLhg1hlrpkBFkgXzooWpR5hAGO6cuiwpvvkyM4dIbTH7jjYtGJ+Mgm75lhNNUxf26fJ5nv4Vzt
RZZQaRZjiJw2gnrFQfjp08668nuYTO/SRb8NleDPa60Y6jkdm2zpVyNN5jceSEytvyvUAWFXQ1di
0iLFynSXHhkdXuCIOPKbDu2/yhpBzZVHnEkzOA/h5nW6+162zv4NodM98Gzj0Sg3uKXDO6tQT3Y5
5US3FCWXBLajcsj26Dx6/daWy46UHwVJXynUCLjNI5V7q/XkJpUfKNI1S9gzQI8sxdOEm0Ic4Za+
8J+k59gcBi9ihHE+RmxNnnDoDpRmUgJCOsoaDWIbEOYmSyqhZ1/hP2zF/XREtBxRXOfWas5LSZhR
HYc1a3HLeDW7rfD9Bw6nCK92OFgZF38AjkfloCf6OC3bvbZ2ZuI/1Pp3gf0Eah2Qgxea1jFGzGWz
DPFkOI55cS8RzCFJZLFj04iVHHdSYGrcNhcFvfPFmklwEUe6f6mlwUCfsUoFw8heAiUz2b9yi6fS
+YbJZI6nm34i8QTK6kkvwVzQQPtVKaPdqF2D47RjAxCuLKq3PHTDhKkIFRwURR/9pm6i2L9C3bZH
LWq6mABaEXn14EWtRRx/nCwulxEWZlmDchabLelMoa4aEYr/AIjJeqz9lUEVKUr/pJi1f+bqB5na
hQRMq7xgCtnUEXHufcmrbkhqp9UOUyKZvsOemDcAQZVqdLSxAhRWthMc8AIn8oLn/vaLKVILvwYp
WR+x4fvDc3277ACCDHJpnyhSp78zfVCN+EowP7KKD9qfKGoSVH03S50JN3hJL8Enzjd7PdgiJ29p
dkuy8CW/bF3wJC7y8mYBZGE4fwrIm98x0OU9hl1dSxdCHdDpSJVw0jFIaUF+1qhYnxBWt/SyIA8q
HV/xpUvpKSOGfi1llB2mnn2q6mZ3X5RG+5gvxX7EkoWwYiplwvtOmnYpwF1CSsG7g4pmOoIIHvjj
maZ6mAeZg8Sb1kQnpbTF+BzXkHccfAGTKeIDoEPmGtSIp5HbBH6vDdWF3vLiejzes/d8PJCJHmaE
gSjACFOl4fcaFPBr4l+eFtsEMaXy7A3OinQzE75QVUm2XxYirK5P+LO1CVYYONc0ylAcwP4SaPpt
dmUxJOiEcmNYUexew6CWXI67bOmYj2WpvRFnEEa6mFPzIbHEZa0Nlu7JmOYqA/qjx7mo2nyuWBzS
BIwa1JqboMZZd2UtoBSRQzY11v0PhrHEZRg4g7AsxmsXuvHyTgiUS43vOyiNbBeau+DQ1Nx9H1G2
yR2X3FA9LkdXeKK9UcOU0papZLsIErzc5U6EfKAIFwrHny9qITIUtv+v+i3Xe7ru1JhqpSHZwQ2W
wVVYHdgbiTkxkp27ZrVXn0vxBX9F0UjMJd9gqrQVHYnKKm18jvM3puDSp9J060rsHX511uI7t/ba
yqc0U+JBXo+V0fcj432rRJr75m8L2A0NLsjuJYsyG8mDl5yMyXM5gk/7guR5jGUPFGzzsBBhh5FB
H6iHFQrV4GXTvDp8Hrq4FQfqYg6zFtgw+xqoqjb2CMY470ZxNe4w065XzviLiZR06EXS8icViGi6
UZ4P8BlAemD6ByXyWc8LOEzaJ25XYiwHaF1IWcYv7lI3Vr0g0YW3hm2sYdxBrLMVBBvUUG2wMAvY
MVWOp7VdyK0ysB3DSbq18OsFMxcLKhJfLIqy9CLdB8YWTjuveBnDafFbnPQgY+OK+Sl0+LxLBnza
bJ+G1jGMSoEIeU6VHTuuWE3pNE4vRzBwbuhKpvjVXVoHgirQlhRpfepDnNnY/2wHit8hXDFD9S+e
TZHFoWww4F771yg9v4neV8RruZn9mE1yghJc1XweQQzjd4wv2h/rRDrDHndTOXslomSzDs3UE+wL
ayX7Dki1hck8ZXMiJKjGveAl0sCKdUGzM8vY/8Fqd/LkDaZsxdlWcD0fXaiMcvP6IAp2QBCQmMrw
H5rlEiMI44Mr1+h+42s5NmROrHoC6u8F4FNpfxCwDgDxX9yId0rhiaXZ82vrFtlm7Ces91Ewajj1
aVD0B9R9L1fNFsInD1YqMPDwc0N+se7V76shD+6mTjGjOY+gIp2LRSHz7whiLekhhOxdaPCF7mcY
QaYHxP2xY71eWWnN0wJ1jkqSitya6eactgbWw2qlrjJT/iw9y7iT1BX2vMoDdg+Lwuu8op8UYKcq
pxsyrrDRmddD+umtZn1xaUDj15jH/1EEU4X+LcNqa9VBO7hDuWH2CpoJi0yC4NFxETZIQjzZkeCu
yH9i1ssXSRxMoujV5HxmQtcyiLNLLF1gRvgKbIQR1NT274uM0ezdLx39bInMqSQqpzOUzeX4T90T
3+LjDEXU/MgVGznnK3lOeG6PobbE+0wFhCPyOZdB5mufBwn3yKxj4jxg9CIvGLLA59lCev930xEz
SzB2zxlQwLeT4TiFeCZzrSeF3gDEQtWb9Nm5ySUOrr7Sy5DiD6Ngz7d1uEhFaxxCvzhaKjpu3XT3
dCPUtTxueZzgHOFmRQ1lyig8lUV7tVeStonf48DYNXsE9aTqML1Q45VBwzOrSIFrXRynopAaqMOT
6Hp8jqFOLk9q6VEv4WwR8ixl/dAXAJi2gOvcZjLqyWQRJAEaxs5TsfKYcuVpWclHxYYNVFuqIXJO
GhoK/L6i6aDdEbb9enmCDUTyySd2GCrYlSi1Sw562vA0DdMFrJZHrFWDJjDXjT93+7nK/sh1KJaq
4Js+KrUxXfelm6MuCNvnY1TyZem9JIMaqD5IcKbxDvwyC+6w4UYLzGX1g1ee+WULZeVO8TGlRBHk
zDtaltxI168q7lwZ1fLBDGKBVza5SracOZrutDb10aP7wzGyIbl7/GDuvEXStDym7/KBo61aR+ey
Jj2dQRMUtuzq1YdUUfv79WSWwS39cwQSWXfbRoyMjmNtku+9+qFn26exj7Db5P38S59oemhW4Hiq
A7Flr2lCd1RhXAaYOzG3PXG9ceI4rEFvDqBZQ0+KuuCsPjwFT7mBPN/hDBmSZC1pSO9CsE52bqpX
6D3sdP2VAp2LwDfAlzYuvmETnVpvN3W4NAgNZwnhSO8vl7lDfrhxWK6YlP0jEJI7mZ4su8wsX9gj
85XPDCaERMPEaiDnjrIpMf64m2UFqaOwvx47ovnaxeVhrLKpeWjc/XGwudYM9mar9HvykQ5QYdXT
ZLajf/CIS/jXe+QyOB32m6Ykn7JWbxn4Pl1gBv6bO6WozO3HWqLiqNUdgkKQyyY9oDlV2JyGUzR2
k4uy7V0l7EYRS5ZTQfDCdTWBjS7tOTGg0v7+p7ikpPSkVfPw6ExpFuWt44w/i/d6Xn5jzcJOnZos
6N+CWy49DCJft9RPclU9vPGSOhyyvzCp9CSyR0jAjf7wEnwskzU+MK5hLnX3mWUyvegiX+zp8HoC
2tUsiRQLwN1aZAaRmHtnUakEo058wz0I2VkY5EZIkPimjrgxKmHMxBjtVBJ0bkei09f2Bl4nzWRz
j4nnY58eKK37XDrlOAx9wxmIn3WQlQ+scAQdyfGaDTNBaglnoKlsEH3MNcjdJ3IF6LKrF3lw5BWo
YP+RzhvwfkgOxekQH7at22k5qX65pfZY8WByPgk5oI5+q2ER+wZBdiygtOA6laZ2efaSKrGNLQT6
YYOfd6sxgtF3G3LDUhn+io4h8WX0lyXp8tuyUN4Jay88aN5/4k1t6ZaJ03Y/qzhhjGnnY6dpJMyF
JpNAvNGNSOqXiRsDmMMBF3EMtizQIlrLS5h2xQAKt8CKtrJH5vYGUx1Rc9R1e2HxMxxubTfXRTS6
8PpVIvJfThKgtHVv8ncCE4IkFYcnb5/kSFJvHCSd4foMQgkclvKYeWYUo6Ht5ZVWeGOBSxTIxgr5
Im29ehoOw9gePD8X2BwKBdHHT0Kn7/lk3AqtjeQU2Os3l7+XuI8V0IOp2m6CUpch0PAAcNzS/b22
QyX6dRaRaQE3iDwCR+Tdwgrk/4wN05i+LDWyOqdxkJSPat/gUlJwWqNvmJVulmtSsvuG35t8P+JO
YtzxAsJ8P6gfWuBLactsojTQzw8LuN2/p7MZDIPCFgNif9oZTnfSvJfbFIf0OEgKZZwyqMhtrowK
5UDCVlpyfRTSvebKQtDGnGMrz9SQTmn6X8pYhkmZgsR+yU/3YNOEZ9BdtoVAZxd9CWG4//Eir/c/
W2cm3ZEgEksaW2+qr4aWd1hVnHkeFwV1tfh0bbwS58Crxe8LLE8dDHBRNtENzZEQ8CQkkRpOAriL
v9j6QrIk3nSQi+ksU+vLr4Hl6zHdH8BtoneYYChdQ6g43tBABpy5vMx9vSpWdJ+lTAxgBEpABdtm
F8HlqkVMovRX7nUdR7MlUXcLZ9oKDi9204hvNmh8QZ1h3TADxKrCi07ZnEN2D+qNh1QwUQzZ6Hew
SWa/BzsOYZ4xm1gyrAARo9slEmgA70oJP82DFDn6dOf9RujxuYhQyISviZrWdyzVuGgSqT3CrJJv
bUHo1ImGpp3KpClyAN6EQ+e8YSFtfi/j5GK3YGIUZFLsNqQQMeNK12dJSlxf338M9O30e0DrFkm+
uqmdg59Fhv4a8hHOkiket/2kYcK53UT4KS2DLthx0YWX65f5o4PuXJdB5NqnKd2fcmwO3DaT/O8K
0KCTGFi6hSuYRNYvNPZAj4V6EbuU4V1c3BqUx93ITcfmtrZxDUVHhAsCfARRvEpVjNp5RZnv1DEt
5hgVzPAxtzAJvPD7PWZIpvrhb4fr3KBqmsRUHQflL1/TxutQ3+IaxXzolHoilnRoLeOE10I+8xCV
0NkqnwThPyjcmtuVAnSsJ5RhVjzkVDNlqJotdxeqmpMR7zBWeLTzWwbtre+KlYZn0vheZzR8zIa1
9bPmlHWQrPeie25kIsZLO760VQ+/SfgdZLxUz1AoDcxxJ9V80Dt54A7SYqAFhRmU+LHhR/4wr6Pq
rp7nOHDomfZHDsy03TwMmO9ONEFwXHCCoxEtDrta0szYnmvuvg7bQwlZDXHmbvjpL4GcRYA2m4U3
+jKHYbl7UInLB50i4SVlR6g5FPEH+hbzETNnJhEvOzi+gJkjTHlARNj+6LAJK7g9OCJ9aQ1i/0pK
4GhCSZuGhOvX78j/TZfDJeEZ1E/TxGYbxme6fQgSuwm9eMd6rJwYZ3wlt6MEzIbAg2phJnFCgfzW
I3DE8XXBGDw31Mspk2uaHbeY45oezDjkWH/eqgtjYrkiKkkfDCENtJKb6pGE+L76wPq00DfvLJcG
wcnVDuEsjspq36n7QDYmuhD4vki57KIvdasvQOJoZi0IS3Xl4izfXgeD+9spuxDlHFnbYiS42VJl
tw6jnTI3rBCQU5zBHXTWY7ovj5Rk5GjZGRs+i74qxr7X6dXDJhpnp7tlyKsXSQxoW52pUKMf/TUE
DBBuioWKeyjmgrJ1ngh9aCdZpzSoAbe40vjOloT/cDlSOXBA5UHQLkXwSCU5IXn9Ry/igX53uUok
ise4A+OyzWwotNUQ/XLBKRYvOKlRiXzbCX5uhEQ8L5dWEUx0zSM92trDr2n6+p8UJGXzyOk1GPzG
w0G3zOyM7/Of306GUrM7n9uroYY/ffJWqpye3BfjtlcWq0RdH3xKvFFaXfRRL4D6//UUN/1bi2+4
fFNGoKaDQdTzy3I2mB3GLq5v5tMcrRhWCEKAkLunu336G/1jA4kzEpwvNHDgg46sv8iNEH2lBBaD
COnD8mbIL1hVE+694N745iF87QYE2CKQKocXR+vOiGe26PWCreznKr0uYYsET4UwNMSnhpxyts/9
8Y9cQkR9EmNf88iVUhOJQnva6TV/r548NBRk6wDyM7VdmPymeARhEJPSyIk932el1P1Jn0i5ZiOV
rabyJ49d6VlcSIMdzinXZR0Itloh7vC1FIHZWccLwiGXDRMxLBhIKE5QcSBtJ4sGXQuBhE7lckQj
7U5WV10jYzIeOnuwct54eWdz/CpWzawm+qsXNDYccBMZao/+KwwtYwZU5CqmOPY8WTHDcvqm1zBm
tWOmn5WkxYRWM4xLlQuLdbrfAoNybmnar3zsEWV6483YsRAL1Ln3o0hTISeYKIrhGdCh9qFx/Wxy
1TDHQJgUsisB4yHubDeJSSyTAQgh77bmEVlhER+HFHNZ/1Eie7iZFxJ96ZBjosJKJQ3t+7QYqPwb
DZP6x0BVE6dE7d3ZoJjqXvtrfh248J6xHgsArtzJWdTgyQhDg/7piiDPxd9xwSoZBGPiw1xDCuZp
BwZevEhCLEE87u3T54+Wg81O0B4f384jBYJdE4nw6qtqAy3hwkB3jHAny3r1P/k8hB/1+0k0+NjZ
Tsdd33Imp830uDkXBrBcaIuO2ALBf5kuBxdvKyD48T8H+qBvhN58VPWAuG2TTf7lowFvDAbsS1e0
Es3UQtH+VirpjM1rGt+rr/zQWyNNsX02nyK92njNc385dd5QnfY92cQVy7IF9NEfMzl1V1mrEEUS
SGdGtUS3ZPTCSsWHawVYKZcaJaQo/D1frqKoTt3LPvQX3yIIsg/qz10HM2cOkYhtVFkCjPTqs4JW
yr5BCrRgGFrk8D7gtyVQwU5gwzG3//lA19cNOwdB2uh9qG0uf25YOHdFu+NDIW7HuxESKuO/YFyO
L/5J6wkiyrgkN/bHRcQ2vIjpiFSjwRs/sD8gImR3Guz7i0rqnLxkh1tFrLJG4aUh3Bkk3teA1ijN
2xU1voK17lSrG9EIEUBLj7Hq6eAIfPceM9ifF455T/7IEInVigvzKrl2a2THTnvyMuwJb60shiwt
7T0MDmDNYehVyf92UXQ40uUJwYDriCESXNCjVFiB2kdw2WWkC209PvMJzDRZ4DFVFZQVI132it+6
q8ule/SK15RUG/+xBYExRNnEHa15QkrLwTQWo2PmcmbowYz+X/LR1+V7t4XJiBH8rcvsaPmb8e4H
mlMGp+YajE+Ps009Xt/IkXvPxr885/J4Aiw46Teg1wuPmvmwQiGtfiseBxDWsP4Z2oYPI9AolKs7
gSN0xnz6pUVwCOaOcns425ILSyJ8Rbq6WaavKw7ie/sKN5wnN36IuYgorEN495SO40JijBG+qjFw
c9lEhzG6Q5myUdnsnv5oygFUkD3hgcaWYZY+Zz17YNPoHF+0X0JyGLUiDqQFyyee9tI3M/Jvk+M5
+4eRgmCd0OxvNhJm0Xu9pWm9XnoKTspACH4EIyZqBVyP9NhgdiHQecpKREw/mLzZCPCzXGsyr63j
5iu9s1W/1NFBn6ggVENpHetSKL0kQWn//8ycGbGzYsBT/GhG3okA7WamQPqOvu/GQvP1fQ9DV+S7
grMDLjC4ol+hu9oxQ5KNfzDM2UuSEKeAMQsRxjjEl7PZIM20sKE+ZLkfa0ws0+q2D0MXpj83TbzL
0MicuP0s8/Qrev90kInoha3nxlnIu8ZROVrvujJZLEG/vSXxg8T5l5wr/zan3LUSLOCBp2wRiIwy
4jb6GVZLRGJfRy09J9dyhQVgGcv5cxLaRLhq6gtoyQuy1b8EIVidAF7l4ndQPoRd+OkgBx/sAqcu
choaIZZu3MCQr0J2KTbBRV9ELEULUNSuhB2hda+D3L6hvk7d1HHS79kn3kUr+BnIaMn1UTS7F2Bm
0DfbB0B61/NACDSJ2CnY1Hx0dIAh22RVw/nSJGxwzo1NLtb26GARHeHSR08BJ+DOdGoFJEucBtE4
8w+tY2nZT/cOchYwFfvfS9sHbizs8lpXDI9V0YK9JmKOn7w/x4DnAFAww0iv/uf1bCjyeIgkPhux
xPRO0+15QdypAHmslBSrqq81WRWt91ElpSmpDlE6xbk/mppNFPrr9Sb8rTpj5lokUS/BP2pShAKh
b/pSNn4Jpw19JeF+Hxeet325/mSGXicxtlTDJa/Sq8xzXFcHbRasWY8MOM8vxVaBOgtbdB1P3QSf
I0JlCNnxCjhUWRsqNPS7o+fM2mZBzgm4rgxOgHs2f2W/gy5LEAB+roFmBsdJ0YkIT3qLfU3yeW8p
ESxjYqS/7bi0nCxLsLjaan3m0gMnVwA7vKefiPYtahnN1f1ZlFjO+9it9PKqKKC/UhYAIcvN0/9M
e9ONQFi6x4+76Q+lsxYs6lnfoBu6f+QCaIYeka41CvzFo+HvKf5/fcJhxZ4ms5xX5XZxf2UOzvG9
edTj+0fCzTBD/giYB6iMkFFVAmo2npg7lboXAP+/45w0r1wOK+yELvoM9pdYqchoKqFHTkQaNzhT
KLTbDwT3GCIK7qhXpQM1PXKzK1sacq0J5LtQZo/ObL7jmL3S7LLB/L63znnGy/fKY39HfpCA6Uug
Etn/gNILz4zQuKejZjrEsuilcRJ8C9GDu0IgssDtNY83SWjUj9iTOBOz4NEfnsuw+lZw5JEEhoaG
9sWyo5pVjUKIF5eiBAHy5JUh59FDS9Lpe0z+rTSBLvMAjWBDVOzsVuG9+iC+XYWF3hR6kEWGvTdE
N2Nxt+7k63P2PR6Q3IuZTpvcFkuqRy85ufqIgGkgH+lJK27zqDm+7z1LU8znXutXcU9xDSXtZ9jh
bv4bBEp2IOD4P+wKuc4zpecB/7aSHgCvb/Re1Fq/0ebjbl8/JeIG/sILvv3e79HsoKa+0UNzr4xU
FqfwOp7GvZqXTgmvUoiqd+9u4ME0bFZqEqiQc8Tdv8aJuiYZOTbKALQ3/XTAI+OKIz+l6U9MOFLT
RvAyOIosOWjQp2AiWgxVU4gA+QJ/vQhoRZT34ARHAExwAWLDxmfm1zAx5lbdVDAIH5AJp3JNcy5U
bRJb6T2DxuHk6w/+0iUQjU3E/0oG7ABRGWRsHb/pfsfxGPf6Rg4O65vTwt4mD7vTgBeFkU7nw027
UJJWt0xN6HjY5MEnq59FtWKmY+uTTg6qIWcvzKDGGyaJH18ANF1GFRYK9kVW5iqJX681Es8mUYnQ
MZ4Ij3QeAXtqvY3pp7EO1ll83+3NHh65JC3LZQhNG9Xk8UCU/Vw85O2BXqRCPy0XicRxucY9U8Hp
o5/92yZZaQN80fBRmOTpOAO0XhbpmyIPn1awdqrEi9NI5zp+9MgOWgI0rbNsviCPEX+/5BHU35Gf
gNfQp0wJI6GWyExxwxMl6adVvQ9/H7kZODeYaRLXzVykn1nGjK6FrJcCc97GS7Ct+1p1j3LjQgYQ
X4KPu7l6pfbks9/D2GrTy/647wO43uxyOLGO7+r+bEbWFf9nilBbVJ3G6p8gVnejvXiJZ63D9WyX
9XGBS1rokl2AAHNepUlzMQj/Xn2zqWkHth43z0EHKcXqnHBWS3C1ok+fw2+YmOLcDl6JxJxQ04Jz
x+0pNA8bHrMafEK6aOVinvQNnIWzTwsodSuKTahR7FLTMTYRMZ/Ew3AjoMGBAo/d7L+oG+c5FhyG
F2dECkor7XOCR3M1vDBIF9Kxom9lG5MuZ4xPGqYArno4HGQsP/rnLWpI37msQB6MmtTd4e2JbIxP
KJNOAM1/vOgdsuq1MxS4wCVDg+JNhCyfvP2CDn3zglkojZ/ZdTKDMo7wovP12jThNmBfyV1vfw8H
K25cabLc2l1Ng7+ZQCMZob5DJUhBdoFTDxUafaRUso9cuwrhNOUkOISFibpzSYqy3aUgLxWt2zdP
qu1JZ9HGF/Fcp82OReYC+J1j+R1oOdfnvCPHJgiqekEj9IwAO7N/s0TwKsfLcljU/G8U4jCD3ype
O1TJYZrmQJooshCmmCDF5ziZyJAxShkb3CFGTa9g6gwb5G/rG1D/CmiGbocNHV8si8SRpSgYu39R
a5bz/30FZWI9uvGRfHt38RDKg3kF48LkPIClqg5wnHW58Lj7QYaNrvHPfnht4EOA5NoGxXmulJ0A
X046+M2TpZp4EstSWgJ5/3bZrbiO7MXv9t//a2oczbequkfsEIuykl7EtagIW9PlxXSf6ScwYzDA
ABEvuCx1blFF3dK0WUMzan1SZUnpXF5pljLPEbd7nf8/hHT66yccm627aiZnR63q75iixtTWTJvx
ckT9jYR85GSMWGWJIewkwcEmJBC0uNGO0E5liPNuKCQT+sxpNJnDWnXMzDVx7ZWZvGTuEw/l036q
OJOR/LW6IB8qLaAIs0C5cRf3dackce5I65jU8oo4dtHq0B8h9fDIXtSgVCxjjQ74CtwcTnvhc9Wf
meD7mwRcg2H4ilpyELGkSzSur2H3KZemGr/6Hau4XMhlnn+D0LGckR6XW8acMVFuTicAnMf/bp5O
cj8MwDc/uR2NOLaNWngiGU04b2Rjcp0vh+d5shmXR3W8Cy+lvuAJPM0krf2JdW+C0HUPxSff3mYd
uH7kVwUawTFBXyVCa3jhoDhCmzeFRHC1268BEO+2gF4V4q0IheQswYWPLrUvMWht10qJp0W7hUw5
d16L5FexgJxi9xRMGIEBfnpTB8HwKF3hselW2HfurC62dPHGePYHT+sJtikx4t7n49Pn7fMkW+lc
baAjK7s13QCIqJbv19tni0AJego5s9enhsX92UK40oS83Snfh6Dr/3Zx9ELu2qA5MaaTOfdO0qqH
WxWas7fwOD1GQEfsukRc6Vero5xtTO1S2qJJYbLfApc1MHiy8pXMz1+f9/rsXUBkn8MI3Tmui85B
QqQ+phbory6K6IAzYSBCceNbYaRCKFgVVgCSSWfCcISr6cLc/4sMekDKLqG0V/xUVGfOh72TpTCH
Ib0zuL0c0YG5EZmgGaxYns2YR2F/2JPv5uTP42cw9Ks0UAOPJ448divr5YV4coX+v3A2ejx9BL+g
O0kk4obfuBkIDOqGi47fMe9VCn9pfORDtuHjuV4TDUb+HyttyE1iF/+suZn0ryDpVT2uT1IdbQOQ
LV8puXnYVhiMDxF/M0lN0fvfCzHVR8I0oZrPk4bSqH9w5FR+NPYQRHtOqtuXd8Dq6mMkbdEaTuMd
850Zl9phkdWhEJGkrA5UCZXvZMv+pmOzs1IAiw/jPDb+c4khvpuvhjJf/H3OGzv09Gz6Zjgt5V/W
Rv3sYBb5A8cEUDY67JxbDweSoGRb4w61J0rQKyqhPlgBgTgdjTdY8ZUp7KyfIZ/51xp72RlnJViI
JXoxIkwfrhtZvf6t9NjS4G7XpShLQO53GV/an7p/Yr3YBbEqHc+2Pa/N9qyVCgHopR8Tx+QnB3lp
20+yw1tIcpIDS7/aXOJHG4CyvF92CpRbCWAE7Pap2+Pmr3FFZz/DbIfnr4Clo+DcD3+VsjKP0d7S
l3Wh7zk9JwRmclbn+nNA3aFKpEG1vg3ZKyB/tjkRRuLkgpy/WycUG40RrR2fTMSH2mnwZHVbKQ+W
DRqUuX+joxH00z3YolGV4zwNoiO5M+rxZxQjASUUYg6Q1KZ3JyME1/1OdOyE2hJ3s3PdVzrZZlOA
e6JORk2abvU+zsFQBD4F/m8WUjf6gXG5PXGvX49Nl5wq83q5sep2p+YA5rCUxbmhSUzpe9abwlz/
X3CwVV+x1dIHYvW+RUO0cm7Zoopc2Fco3+wd03kYg8ZrtiLJCv5lGTIEqZTaCPxcRztxatUtHlC4
r2HLtfUT2CLPi/LPShYpQ1OOGqiUwOS/ysGgJE7TczyYrcbxjP4oxanY7fZPp70NfkKNSaz1QiGh
2nIdIvm8X4IWgtledHcR1BrUm3J+ICXJ4MqcAA4fi2GKJ0upEE1DGXO2BcuVjVzeXbzS+Q/fN0LQ
LbKt/LMKfd3tBE9kw9keEW5dxjgFEOBLu9GdTXB7ms5w1WvmzMXmtD3tmlS72z9CkYSxgMmlTTYQ
9D3J821HDXasB9KfiGibHdu2L42ia3g+UIrpk6BJ4633y6tqA7PshHCJ9G7mQFpMwIeqGXh8olfY
hOsnPCrXGg2mUmzNKmEkMghwNtQQNaxrUmahBvVSPhGzvISB2L8vkpBGgXXTkPTQAT1lONmkRToR
tGNle2U+ZH4wAbPuHCT4I2dNBguYGfu72ZHJWP0T1I2X4n75LTUkZJduteSz2jDWpkjIOL22fwg1
Wyf0usEO4UbVTf/6bWVVAYgyODAQZWvHBePxjMx4DZo73UwCHQaofxSvJ2K6hG9M1zTBbxScxOvL
6e8YHiKBYtmCbsGEAeyr18XTC0VFvm7NKkhJA5Cc2LByk7XrD0QX+EX/AzjYUEZBxVBEqs3f3Arb
QCiaJWYki8m5C+b4tpXRXPBvIPylEOejtJpyd+XmkhU/tNgIOQAHBsFD8twdbna89W1t/w/u9tK8
/VzfXSSleWjUrPmZt7csN92XaVCW/YA9v4q/36Grub6bC4LXV7/msz3mVr6l/9c/E2sIS3KxQ9Qw
FsAfdw3RtXxktB9QZF+UKIQKh/vSSyMocphTEcRO7R0AozOm/pTav1ePK0GqBwOA9AqkFuBWKp2K
5S1DszV0Ms6ubS3btctIs9w2isSvii8XNGHTahuyJhaeSmvPMGcPN+Qoo1yEHMmom0Sq9J8HNbGF
Y8MuBnoCU9wknwkBE3KkEc1R93zqfIJUSaje3Up6XZXslWtwqxWPcvvd2UPn3yN7RbAQjAmUOb0o
QANHeDV3nlvG8UAhu7rLv8tg6Zmr9aI5a8ojibUC1mzL2nWIX+G3r/znNY54fOGLoEEM6gL6VZ1B
cjAyloVS2gESeq5RXdh0JtvFRxSFZRcYurhKGNeR0gRb0FfBvirecSLPwdcK1qv6oAuN1NiR7Etm
N1C4VUM11yIiowutXEobNRrAWFRggKafgM3l+ULLxDnmRwZVx1ZaA5J84PRw6GXznUXZS+Nk//bI
lODp292O4h/KYZu4FPe1Dk8RtNvn29BFl7EUwXCadAI8ePBiJsTzZpnGyPdpJss3g7J8fu/vFF+Q
BdPGgFrtL9eSsK5HIoj0GNEjKMWCT2XTC12ccHasg4igAgNPkUplMVkF3AvJHNW3nC8BksvD6F0R
tPnp/lNEUY9o0ZPt8KnAaNnsNYt+a9Hn3ywA+jiOSih6sMDy76NqozOLcE0U0290q6DkobkrUOZR
lr2YH9ZUNAsiCMKJV5mc2yP+mz0tfjC7e+zdDO9HKfST884pZCahScZiyXvdjZnWaRNNviCcIRoW
2deHBCrjKdiei5mYqcn++MIHknkPY7RE6OUwEnUS+sH8NzK5R3sK1yy5smbYdTpRhB5wtJB3qyWw
NetkyFz/X4Exd4DXIG/+vbJQNQ6V+T2zEfb2Z3Hp7cjqx/q6FreW456/D2rzi7FXFAKxJdTB0EU7
6IEnXY/8vOavuw7ERNXaESQyTYbLwhiPDINMGS1VkEX8ukWxwvjHpl5YYs8wKsqM0Rg5l5A31x62
ZuCdMBcz4sp2ZAKRJUWQ+ieHqLfFlyQ3mZtLg3PzQr+OcXUDvK4vvWP+WisaqtR3Yf5MUpGpMveo
hOxEd7vlxXRd/bu4CpbrUTA4q08FtAoJfl4Mr5yvlNhJvlKOeKTZVchwYwaZ/Jv74Cn2QqMnJ29b
tnQ4lsh3Ck8p8NVUuUSF2FroMbanV4YJ+X6SWd2z8gONmI5MahmI4LwwIqwMoOzJKEAB9UaXhlOk
BPmYmtrITobtj1Eaq3SU3C9zP9EtiTZfB0Fpw9UOJOUWc4MB4If81a4XdY2nOWgwEwvj9sEL8lPS
PKI9/HYka4I5gpEs6ljKRyCS97GZSVuQlz7OBfRhZrH8OZ8yYdv8PrxlxQzouKn41Kc7MQb9IIit
kHst4Yx0AM2uydu96mniFMxz6r1cHnqnAzJJt2eoE91MlTiSfiO6Jvr1in7tie2VAejQvyudWO4v
3SaR5SE3/l0jfnZW9HONhAtqitx79DmWgCn5+78BTHLZvwwfIl+N/pj7ADEGMEGVjVoIZ30TT/bk
b3AQHf04v5breyDfLuPpji7l/2o6uCm9cK4fs32Yl5t6LBgxus4/9WAn3TWyn1Ay0jt2SN9qsabQ
kl5nG80Zhg5f80JXOK/onteEEV2CI/dM846kL6h0o6Y4n690/+YhLn6/tW7DboL/MAaJSbAYR/78
ur+nAnKY/6z+HeOlBCvUfcLjjMs+toW2Dfy0hwqOS81JtqLXNYJJ0YnuAzSJ31+F3449IQmeaDs+
YM8MOqYsRZXDpazn7D81NCq0lWre60lTY8exM1wAsan9P+ABgjtV94WqmA25J3LwLHYCIiKfc5wY
dGFSXyVTn+r7bLDpJ+qTMOrHutgVW9WlY2a69JvExgFRBaRrT8MJbxm+ArKsMmojUDZ0v9EOBf5U
IAA+kg7VL1m1ev3ZLA+ArB9lao4Q6lgmvcNBghvBCvgAfJwKWgYIpZW0foybM5+5RsXECjhr0eIa
dkzixEnWHWDRbiw2NlIoeBx0CgRPNLfggrJRJ90QnWC8AFi8BQvWNGQVFWI5J5Urxb+sYOc2luxa
066wCVDKM2SFaS+xfuX05ssnDYpTs1UZ8JPakFng0/eEN7Jr3MmM2edgVLaFFttdZOHBf2K+lH9I
o7lOXodkWaoX6thx/vb6ZgzCEBVWUJpYNSSWfZyle/HdIgpfp7x0EmyKhNj30kpqRTl3Cfnqa9xI
znMPLIWp9OfTPKLLsZHsNfPSjx0vc4eILBiWw198GgykaaIBnth4qeJ9rzjytYQjXinU5SbImVZV
9tyMKVpgpfOSqou66ry9UwlJGbLyidxIhXoHEWslkg9xvKlsaeYlj4PdxOZsFgQK0zmB97qY0Z2x
+4PSlrQJK9JtTmokS4T11GRezuEn4TQJkQluTccax9hib6zYe7/frutO7jNdf15KWEIDZ1gi1l+j
oJKZfsRMA5Q0bw/NgyptLjdhOV7Rq3Im+F14aVkj5Tx98o/DOY4XX+EdcIB7AJz7BF5eaU6RtqHB
K2bjhiVY+T6M59G25NCsMr4sTabUrGKzhunXNdvOz786G3XWAMtiknad7mT3/LXJOCD02A/5UvFz
35pw2UdwQZfySj06AedPxU6IR3DxE8OozcG6j7U5u1maeWlOsgX8ScC3LaOjCrdQWGAsHApmqSuy
mY9l9rKRSbEO9WO24ozIQvpXaKBnoQ0hElnJHKHxFmvuX8WVXUVYIK18ScwxMd6vNOgXH4WHP4I4
gzeptupaexx5AMVU839YeoCZP5bZuCDwFTjkAu1BSBd8OWubl1UdE2g3w43sde3C4oW6BkPnE78Z
To5hSgrXXCGVlUBVqXROatFASshyU7L6S4Jb9Z+Ucbfs9G+D44Ybwje4CkXWqLE9IJDj3uCph1ce
YGbKz7Xi6FOjcxkK+41kVLMiKERv+hYZG1OiYqsdpSw+nKv2F2CRC5JknotDyRWGm1YxBIzibBJG
MjQlMyJUZawjpH2V6ToyDVh9HQcf101IGKT19cf5EbfeAcTjilaUVIKbs63d1jfLmTHZLO5wGnPm
GmOV41m10HdXeFDK+DMlTrHGeuunhsz6EFKRvW85rgm1ZhVD/bmbsjp9Rf7NxrHD2s3UTYRZwA97
5rnlikv/+qhGZmRyUUVAQ1afNKgVjqyvmoDo+cB2LGdnEfoPFzsuDKbFHQipHKqA0jfJhFzQfDtd
LZRhzvx6bRm/YEijIGMfhawqg3zU9wtHcmf2Ojn+JTO7leFqlzmAgxEOovQ1iqNIkbCB7TB2Sqqm
UDUwWEqmmI41zxU9uRQTsRLJ4kfAxgOXY7OKL9aTCLqjeNbmtS8mnZp4kbDXk81iAyP7uqgGCxDz
SlCfWRMDu8z4LZZ85em6bZ9w1KtVdiwgfOBolGSuTCLQu9BCwfbA40+pROzYDO1Zgz++yhzW0QAo
UDDYMqkpvJs7t6uDAH0GRBFspxprgsHYI0ev2HXfIBag63OZpA3WIQ+XL+CS9YnbJTX6b6FzMHUB
6inVmZPT1ZvyH3zNvTdDoziBcXEQptKNeoaEi/9oGkKCk/7w2lXMFIKG4InW5NMX40Lq2GIehJ5n
jj7H4ILKVoNGcOuK9emcAmIuhE5tM37j4RVmFc/VX3SbLyqKT1OM7lL3q+BN/z69gXCrcRwoos0y
fY/lByUca+jlAU4iJFXduHrZX5/Pzg5aZVWITWhv+t/lTdiyS1mkE6v3V1QspLAHYhJ2dARWPQxy
w4ADoHChiyNzPbqypYVI8X/0QW/O1gt6czT6JDYAp1tsFdD05O0CostGVUm5O7XMgFUuIF2N0/nE
nDdPa/h9kKUdfkjxXoDgtBFSb1KnRCCu0VpTOixnue3HSUErmYQy+wt/l4QwNDyyHVq+5jbWlVeG
0G1fKPm9Z+nRZcg3FRVZvTkR+ELYndaZOHP9ajgI7sYG4wmlHWrTQhfaaRkta9OycD9+Isn39Kgh
UYXx5GjL9VdahSsd/sKo90jCfMkdfd+aPPcByJ57jATM6y0F9r2KLtkZAKAq7hsTDqgdts5YAGxJ
rvCPuTt5Tv+IyaWunl73DwWdtGoBcatFiZp8/wouAw8lZoeCyxIJIEDCAxZKQGU1Hmga09kXsUgE
7Q61FPu6um9yaCRB+Q85yKajFNCTnJCsslebgaStb4xa53cXaRhxICU0az7QSXN9bV6CNiSBuPky
b46tOvGBqKyI/05Z1sJyU6ADVktSU+iz7GuTr0oXZUJ6ZDQ6VHMyOb8TDp6VMvAhLlmLgV7zwAPy
nFaq+xbl5nEB0eAn52mbenlhNxN3eHOjYNfq1k+11lX0uwI5Kl4ugK93k9TP4jG9A0iIJAauMyvQ
+Eux2s1aQyOcxtXIXkHZKfJNffwIPYPbPs5kPlpsLhjzzT30ZyTNKzjBGQ5BdNVx7IkNjfyvETrm
v1ypH0wyo8MLnZIonziFNi1fJb+Z2i50TD1WnzDtoL6iPCa0dYqjs5RQQKu+ZW05MMUVwvD+Kr9F
XmcqyZZ0pfdvpM1GO3hRBUhBUNdIJ/cAnCglco3TV2rkd4ORyF0ptMH3ntLBwMtopcbuBtS+KssZ
TqROwQ4BctVrv+OZnpuoXS1Lv1rGW9CzmvdBlG83FAiAM96ac0+cjJpfA5u309CxvfjlYx0iPZRU
gPmgIz1zEcwXalGi2pVAvm/Rva06JZ5tTfyMIEqJWsZP4wsO+IYFqfbfpsWlofc/LnOuLTaZNZ6q
tTLdFKhJVdtCnck1ghscsxWNe4OcIjbW8xGeoJdq9dLisUmNUtcHQNCdgA7XHfquEBCoDmc5WeUG
YRgtD3Fpb/AEVBeT5tK3bSCK/nka9YoO+TitKqLduLshTcNAYsmE92TiTQ4IOOa76LkbMtKvtf3Z
Yxkwke8hV4R1UWMKuKebGrewkzbhagt31LNLEwoHPoE9boAsXHO7nLirHmah3ILOHOAe62ABU12y
dGozgY5S2GgNtvKbmZoNzb9xMw5EP9pOTnnsUMR/mAGxbonjMpH09i9Q9984d+lT6WLPgfh/wiCW
yuiavPPiHMVshFYfhCuAJ8wNgp1VKvQUN5wxsbg48tsFiJaOJsbnlcIThsnVur4EEnSstTzkQevk
AqpkkokbohygVSYQ2b16rkexzWyOKLuamvNi9qP3V079xiPhA8nErHiv9x0h8rtiTlbTgBXGol4B
sXem7NNyMwca28Bz/rGlbJRHN8o3rZ+bKry6RfEj6g92ugmn+6QR9BqParqwtny/NrWkP03kQXBB
kxWGDragD7mDbq2FwbBPXl4zt1rwNb7MLl7kK9/lUq4X87XXPUAlHL/iZuvRsL6wQFlWEMfIHwBm
XYJBQ6Vb8gdYWupHRWpd2bUdJdcH2f9kev0DJ563uMTDkMZxOX67kAjLmJsi8idk2w4CgAYEE/ic
yTQ6O6p+zpv+5Tyhq4TlwJwPj6AXC1tpVnUD2JxI4uinjwVHy8JOd3JKLaqgrHEJBsMr15Bzvt8N
aOvsPaoZqIGJ7sfjiTooFr/pKnDhx+z86H20EK8XocsKytr6VZ1CcHAooVDV5NGfKINr0iKXBpgZ
+lUdYKCH/p9zczRYwSXJxwezMJBFroj0wEJclm+TWvVrMiyy2UQsvW8B663rlKlXIIi8lcIwJCdU
ITa1WS4+ZiZgovzVNl52KBf9JbtTlMh6J/z+ILAH7GFeTFKhjzh7hcPMs++yEGCSEZa+keEyB9Ui
++Zt3wOV/jqx7wPmMuC4R0FMFeMtWYKVqZ0oOHm89mjND7I0FfQuZAtX6vnhEYiVDFbRQApbGO/j
pgKhiJbghp4fOOJCAPMtFd3tbaMkGwxbFhCFnvUK67QaamZcOnsh7VA06Bya0Vy0t78Mo0opj7Sq
XPTZO5Myvq3QNxstMWQzIuErR14OOeUJa8DLto4VV7mibK+24PCwscd1X45I9JnT9peh3DkssmQw
t9vWKI806/lkft5dsQlLo5ZOJ31vNhEI+VbSIuQp/SLnmqM6qbuYYKPb3UE6Yxf/UZKRMt+Zz63h
z3PjCva2Mx9Ict+emjdf+1/0DTisPwxRX7nw2s50qCszw9a8xvWuFwRyreSIupNP/LoqWa6sYBou
Oi7gRJW9jG2zy06upJktoXlMiNNjJw09FIKRROvW2eoBAsuLkV11yMr3TOwA2uL3LPKjqT6tnDA9
LOOClJLovtvT2BYpntkPAvtsKpC2byh706oC81+KYfJckcfQGaVvV3nXd0zGubF/XdiF0Jxzc4zL
890tLD4zoUzSIFPXwcuSNU+66ayTrNs5Eo667jBEEF7ApT3/HfRs4BXwTG0gC/4gnb1vlbTWTq0O
qTfRq/ImXA1hAjTwBWmcLwFGc9au1ObtPuIDusEKTifpb1hcO2JpiVFd4eLgdwRjt3aPWR7a7J23
9AREOC8/kQRB1oG8kwHlEBa7aST4UV8TtAZqWeqfBz91g1os0WXQ9xSpbuulxaNzQyWKYuNWd/Oo
b7sooz88jTbwAXdQJDbUTpuF41v/1RoRIC+Qs95ufBmQDIGAgCimY16ac+UK1nJelorfZFH5Hnb7
r99rL9pa72iJosPyfg9E7jJwID6RawHZV9gbhvBJX0kJwoO2CFOrr81CE0n4AT6l93GYaykmAUZI
ugyq6AsqSCfcY2PTfCi45XjG9l1jfOVFzwVGGDkxjZZwMHaiSiTfMjSAiweyeXL/6jNVT1+ljyqo
h1ODWPNZNQaGW1zdFinktgHirbc2XpkGidLyenYPIFTHK/7k8QAH+3LXJ1CD3g529ESCIfDtecI8
uqeNI3RLKTSOlyc9yNsmi2STd+9OeDoPqlafrV/K5xxEFR9zAuPYyvw1i/ndOA2XvzHaPsLAY9G7
8mPr2hEj+vcUVLe1P9TESQNaJIspnrw9O29JbOTUy4fRcqYs73KAUsfQ64ktzBhl8IrQWI4Jr9Ng
GwMaG/XGyJPs2hdYjVqXGLk0VY5BYNuGx0JnyRW1f4EBy3+RKD5ngA201e8+O9QUnk3ic1vmVwC+
n4XVRaR4BVIDdGxRj1QPTomG1BD7aG+Z7cC8njFrD/LW9LcdUVKIltc3Kc9s5loBhIOJCuju1DSX
105Y8cu1MDIPUDICiIWeo6sLWRpyQPd1TsEWkZjQTbmWngmkva42PN4WZmtR3tIY/it1f0I8fZ0X
tnTIppHVnSPM385aJh1mWsIGzLQhsG2SgYzgdukUWqmU4XChIVbxY44RUuckSO9SbNWBVW6AlvLK
q22UVwPQb9+LtBbrLW+9IYoGlev1YNHJVwctZ57uGaUmYLpseEuPXzEEH3/WoBnRSWIvvN9nVWv/
RhfrEFsyuDPi7AnyhpRBBbeEiHTp6GQ0LCn8UCCcd97aUH5rOrP83bnHe9WTSuCgqd1Wc8XFPgSL
wBrRxQALUWQmE376FF+Qrhq7i7agW4k8dhAPCyx4tCatlDozVQRp6Hq+DHDolCbLntTRMaSQC759
Mg0y97noIoTbsS0vzQBOPDNdNmeiZN0GtnaaG9Dt1249HB0zODlg3NdmqnbZ7U+86L5YfKfS8yRS
ANtzh4IqOTDgpBFBqj+Mt7CZUKM37A5E+Qvxp7yP/UUtMMyMpXRBR90CmYg4G3svwWszNyt5AdYW
/BM25EawwX1IZL4NhiGv5R26ROJOBhPJwUWuGFQYdkAG0PwdYy2Hj8LRR+d6hTixBlEVYy9cxeEz
eWVdwupHjnXcVzFtJtTos5Ne+9uIfyswpZ8GW5988hIh81fZArP8l/pCVeZBKs9GJPRdH8oyoRyX
9eeVNNkfRzrCzYpCwMhNg7jYvaIIc8jcOjmlEx6ISDBehGpJxiUoijaqSaM0Zteb65YWHXQMNR/b
PurMNy22vHfOLeBrS5nNTve8Ev9gwX/S/L6n2N1Cw53cpUjvtBySNag2NR0dyIBvOj9N80viD6+z
Xw7u4RNPQWn3f19eKfIE7YZdRcZhVg45uFcwmsq4o2Gb0sbpqBD+ED/hOl7IKjQpBc5RjGsEQPt2
+QoSpWn1VFlU52H+RUNFSa7C6PIBTdSsUfQrB3PZIoaSUSSEPOqQbaUsYqv9Q+4wwBs6pnNMWGYE
KJiFd3PVlVgz5hks1TozyqNG5sfoyRt7PNVjwrFqQW1fhP07xxKh4vDT4t71TZpPY63JJb3lnR9U
dsOjGKL6iUZcOT6jZNj+TY7W8ZPpOPu0ykTyKMUnU9v2fdyUVBhCpy3sSAHie9wQnFIkQZfrRtBD
8FwFYsQc9W3hvVCVvq18pzf8oj7tNLp3hS463SEb8aRBfBJxCG00r8sipm39t+pA3NcsKC+E57aV
bv2noKoeQE/jT/8KYRcpkggm2Bfv4Z8Tq8BliQDdmaWlBBSF1WUAAww11cdtDtMIahENpQH6koWj
DZkMAPVCebK6ywISzfxkfENkWzzRD0AMiYzpskI50E/jlwZUeCIC74Iss+3/6HHJ66CGecuJi2Cx
rznYLc88+bvldqAF2uKxci6Y4z8ryuYFFxdfeivGftd8Eh0AaUmxzI20PQEOXpbfVZ122LAIQF52
QZkgkEGcWdFLN9xO4u0ZNlALq+6hpPqJxgzwtFFnJ6X83WO/0P6w8ez88rjGbQBx+/ihzaoYQJRn
w1RK1jKYwPyXTRIHMd0XEUP4ETMhWtgDj6orb33W7ILRkMtnHnNVPSiNTqIkthAk/+dCY9bEKNeQ
jL6lNR20FvsSWLs6M9Eqv9DnD1zliUkqBwqJ5Pra8W3unqCagDYGr1s72kHuAcy69nkmlrjjj7Lh
I/Buf/KS2l0vlTstcutJjvvGJGjeYZjqzfKJ2Hf789efm2T2RQQkZ3HSe1iTLSXIOY9QmY9D3dYe
+Yz/Ggpkb1A9uZgk6Gfa9EOwXhTbMe0NxhfHsZwjEbsNW/M+59pqE6Wv6o8HOxTVouhfIvPEWFSv
4UTHj70MNByxDuqyzaOV6TTS28E/PJaW4yLXdZPoGKWRndGUzLbHQaC+jTq88QADwjEJXzvky1mi
x08M4eC+PY6RewN3pqX1b5Hp9uHHQ4JgzN9W7wVDQ1Lr3R9/5N7NyeRNAr8c+PGSOKXsBjAsgc6q
G6UpNk15DjckrsbOMyEI++ZSjqE5jvXvNETip9NxRdejtvFp0chSUscneRxQz5J6J0YgerXZMR0U
ymZlHJh2Vksal40Qg9JTF1V0XpgtFFW4SyypLEf0z+jdJhHVkrzx9gye6VL5FbeOK+cnZUZuHPvJ
eOUek/aDHwtJzgNs0YiyLkaVtGT7oSajLGaRoiiR5QwB62UUbYyi2UJwJGzPt6rb4iB0lB13p9nY
muNoNeSncc03btHFWZDiLEXAIdainvF2v458FqybYyQQ/Ijsn8YaAvi7LxbOgbV6OlGoJVC0k1lh
+nQBOKOJTLszs6+ml4uc+ji8++Z4WlAlk9F3aBtsdVaoOXONVjJz+ywqRdjPjMYVh7sQJckUC0g8
V8n80WwpWRc6KzA02TCRPJgMpMsmQHyLCXZhMRX6mnI0fEGmlOvIjRB5NaFKKvEpvH1hLg+TY3WS
08e+1rn1RkcBTnmtPLELRgi+9ybMf0gmaTnm2Xbp/1/hcCOJMGg79OsiWa5Rzw8tf+S1QI978PBv
JBGojigA7MzE6ROZHJL+cTX/73+STEyh+g94bXSyoNgNUstshRfyC9T95fkCK10nksmXCRnxFhUB
xjVagxM8LMGtGjExCtBrzDwg1wmIQL4icSwz2/w17qrUcd7d3FXkUY72ldy81ZctKhdNRrg/Xi+S
2X8EVGj8J2FtMpC41gaHyROi3IZECtcBb+WSbTPzK35Lr1j5Qf9MI/HNWCIAHAKeI/JYcGRCHpZB
2jKVvZwxmRp84McN8ll5VYSqqrujVv1JNu8FU/Z59bSwbsgGBqfZh4rQa8dbU22EAbKwfBry30Yv
2Se+9qeaWVv+nEoCj/Qvr7QOX4xNa33jSTNMAFqOcPES1yA8F7mppquktlAntKRXK3eDIO6IC/HC
6PR7Z6GiEQBD0Z/LZyN/6oCxom2mklPW1GnMx5ym72ihNI0sbYUD4J9CTQGAb0RQ3cszk/hNgCFk
N4yU2gcrIkvGxVraA1XxtNK4pQjTEq+X3a+NAibmYwwVH8NocRNqKstjwxN/0OPs/czzwuZX/Gu9
83qAAACWQba8vukqCrxXNI7m+cQETIn8x9I13uoztCpYvpm4GBZ75TQtITA/Z7OxmA7TcvL4FP00
6q/qPaMX06Yh7Yr5XWT4KSE0K+VkHVLy9lkXuLkOPPb0XDlcKp2xpKafmRJr9PmAbWpKgJYIkFPe
+rjmarc46b2p7tQRCIiJtqybrEKi/kQ0KMP/Pjbnd7dJLtpr/njkgoD4qvjKb5kzPrKPBwJw5Pj8
r9/FOv86c/GvudGUbt09MJ3mPgu7puxU5SVwK5axX3pSRXm34zxKFNu7UQ7T59mTlwqe2RWeX1lU
Ufh5X8hYuigBRHMOSnDNbZtqtKgGSPbjICfeYjeMWJaXsx59SJPTc9uRC+nJyuE1Vq5WlTyOy+L8
HQMdTiiSyMO+ARGb/CuISv8vZpYZ5G9c+wiEhLGmHM3VrBG0Mt/A7nYeid84OAAYsHta1huayfqQ
idKvtRu4Kgzl4skS4khmw1SnAJVRE5cj9bCZPR9oJIjGo2T6hiMFvq02TdHnUp6/CSJvfJlMdr4/
WNBWaN4HZhfFr4jGjFoCUdccf6yqkf995Y/ewvaDpjXQxQa1s03337zAs/U6C7TmN8vgcH0VTPIW
7E6E/OXRrzgza4Wgkva2EhpdbXi0k3MN2sV+rY872lqFq5NbP4Wg9nc4YYKZXxHDz27q2f+AK3lQ
OLZChyPIHcsnqfeVwb6vbYEksPEu5tif9hj1vbfacx3xzDYCeBRQ7Eg5gBVtPyhaKfT8RkBDIHf9
vJ4wg5BGRipSEpNnZfBSQVpfS3bkApfIWxiLF+5A0k6zRLR2sB1XNAKYnd6YfTUE7f7Oc6fmDJMZ
aRWwwrsE6glTqQFvCcl3H9kpjmBLzlbtqF+fK4IBZ/9/XctSL9ifw0aNZ9qeUgw/berIYGv5tViB
8fhvzpF/nADaV0cpWVlHJllba50SDmA6jwsBh2GtPUWL4n+3A4ZGWxy3R0yZ/N/Yw1mAzKvbjE4J
+W7xtwwkCZgNGXAAjo8ZnLZZ3/qb7+GMsalJSqBFNjaF9b4C34oAGDnPDiY4In7O6mJ/r7ETIPco
i+TL8KkQlEjvvzmiNptdp6S9kHInhR/6nLmCd49bax9jkcMtl5zsVqRW4J9+dBOuFsCdE2FDMoA4
XaUib0SD9z03toTU66xMZT8NE/47dHsFobSwlahdWhLrRb5yYSGoVQacqGPIQ87HIiLnNx1cCXUd
YoCCoC2fJ8fIefDFLWTXk6S+f68DBbCtR5osvUljrnpWBIOLlt00j8xtGLNOjfKRQXe6f+6JCF5a
la9xRsx9RMS24wqSoXiuXJ0dzDHDYcA5nr6IEktQDjZelbV6Kmvx87zG+SALJaOEP8EtDjb/QSKz
Tq21aLphlG1+NRR8SE5oKSbOb9EILWNaefcEkNfnQpS+mWLkrB69Kggutkzt9N19Xv/eFYuSn9uJ
DgzzmA2UpOASyjyULVCqF5dcElyF4Q7vCZf5Ifd+p6Pa+/onFAKy5AyGKEDxQlGxfzwIb/hEUtOV
gS06wPK0naGFM6BEZh105BYMFWW1xVl4QDM41E0csYcwrV54plbx/K/tLCed1e2UzUCZS/ExFrFW
oTfvp1qz6z5gwyqvdcRdKztbekSXCP0vGL45vd2d0evA1x9KXp5xXkFMqpHYg8CBU4IrG3JAfP9f
tkZppgmugJYCgUeusFdQ7uZFNaVyxbUNvSGU0fpMoCAnZTJyQR/TuEZBrBnAxmBt3nbXZuwcn1j5
bSVL+eOvSulOQUbX1Z5QjjqbrVzsFSWtQ31v2AGRPNpRKJHAtB+QtbtrEVaPMAPRGNDY272TTvyI
xt0OzdRkVPvUHGccv0O10JTAni+Om0J3NWNrW1xg37zP8g5Z+GyB+WBJsZEM/bNQ07IrhZSBMgc8
mwZ/TzNReW+UKltSPPuNE1TRcMwvDuDf/t50lYZjp9VBmP6Jp/oVSjq584n8O8w2IJMOgUu3BuZc
7v15ZnsTZ1Y70BsZRC8xakkWx6sWwA5ytZ3fVlwCiErUSP0wp+6PvSAkK5w/oRyClJX4K3Fnm2Cb
v2sUuT6UCJ8ng/mTMP10qV3DG/+mD//swNpe1IKBQE5otUGywGFLw9GWJ0vnblci/+TjMgNaUNZQ
53eixsZbJlWFmYp/T29WF9PRJBzfNeZrMH6GdjL+trhFdHYnD91cVGHKbuhlmRtj1t9Gtv9qdWko
cRtUyCJtgJGjIakUnEu/L2BOfQsGfdMUpVPF8un+wDLzcbbpDZMUylTsWN532Rgy4JvOL2TpXFzC
QPw1+fSqtddE2T6K5R9BRNF26qXASeJXhuORDy2Woje4dFIDLL0iuibFd+cEa5KqNBI1Nx0VdUTM
3SwV7Rcxfq4uiDqeUOMf16s3D80c25LpdL/x0ULxH18nQ+PrR1PbQ2FIFQn2K07AVIrg155p/s9o
Pg7gp+w580KG329h/77AY3KfwNy4Lk+pThlH136VZXucKqZJQyT0kkUsNGqE+EVzOuMoS7fxnZ+s
SZEQ+eyxBiDB0poPCNSms9KD5zQaUA71mGQpy/zH+Z4u5fJyJeRk3Uj0MzlltAGK1QRR9CHSMPvC
aYyCjjSAYlBerFNskHyDak9/0jc3YO6vZm1c3NVN1ZRC9SIO2AhGM+OE5IVpK5VLLtQ8vIa5EJS9
5Vap+J3JavQDW2N4yjPKOIltoQiZvTYmgKaRhlO99p+4EmqISxJ8x3jCHNq9BlzigIu/KOlODGKx
FBm8yhB1Z3RdGaWffPUJEb1upUUAd9JRrdyZrGenlF7yacVDGSge/GthAzBa/pehkcTVOAUIswYz
tXiiydwpr+9vmce0npJ3/gai5dMSFq6Vp1t5Xh+wzE0V5e+Ha8nKA0O89DWQJVsmhw84i/+o5a4R
ACVOQy6MLvRcQqVeyQW3M3wSlg0sea+qYuFJnKZHFsJAh6W4PeB4kCrVlyrIkUI98LdC4hsqceYy
/9bplJTby6ESNKPNR431fOeg+RNTuQvh8sKNIVxNdyqamCqzm0Vptm9HprmhoZkmDI7vXCgPv2jr
tyoGboLFuRrfWJQ5kPatVXWHaMySXqowqf06Xmnjc4p08dUZ5hsVOoRKJivQ/1qP9zXxgYm6/a7P
NqxBH/gl6sBuEJ8ZI/PjblZmeBGa5rib+xoMvoFD2ryUVY9KfbMHGiDi1S9MKQOV9b5KEZuuxsUf
cQDRpIBGJh5PLZe4C6McHuFxHpNm772wd86xZSFfMvV3fU2U9eU2eM3XZczwLiGcQPu7PFm7hvn6
agypeGVgCfQkHapPyAcjeTWWi8Fvs7yE7FOe3uH7zaJpp8Vr3/Ei3PDf9d/CIc8PljwUiTGQwBvp
5vBLIEfiaGO1O5zin2nT32u2L/2d0OrV/gqB5wbZ2akvLKlxL8/NjYTpPudk7Hg5C2CdYd43UGDp
TLqOLaDByG2czrKDm9OvMORGGY0WLGsaanJ4codvdMnR6KNJe8H+8G3d6TCrTDOp5vvsa7YlpbV9
Gm3LcyxXuyyRCNxd4YcO30IdLOe/L5mj3LbR7xkmHhMHCc7A0AQZfqYOge+aQJnAriiNfgbbljax
iAiLc6SuElgD+Qust6qF3ldy45ShDUJG5VxuuO0RaIjC4iS3um7bmlu+gIAfsWa928d0uxTX1Oqh
cYoYZ/BYn4ZHGW8WhFGLNCub4NW9NXDubA/3DdIj72ZmZRplPHLci59rGgcgVeKg9xqB3iLCn691
VCGlFiagEBcor4TGLBI/CSvkO/cJE5GVNsAv0ZrbGlVksjSjODyeEGCws+XvQmkWs+o9XkQcWI6M
tpRLJ9HZe+ZRYn/scEIV6hCImylnO2zuE8qx/DEqocTs9cY56f4+IX/h26nC6zPm42BOblUz/MS9
+QFv9aRqjBgPF72SbsiB1unZAJer3djRREVs4/VglxUbgkHotxo0ZMDoss+5YoxXR7CtClr8FS5Z
OWvB9WAn7KWyt4LDHV9DkttA3A9AK9rncvqgYjcxG634WGOD0ApOfMGxght93eaWTd1wBpDDbe7u
jTEPdpH7UUvANqgzAbF/otUKiZElM+U3sJjGNv5r1DETTw1PcRv2vKBWZ+DdZEh95QNpmY48rEHN
XbtdsGMQbghXEMzrL4l89tpxqdiEgnfmTUWq3vqMHF8aMcivMOZW2ei2y6vAQ90mnTcdGzQqOiDj
q/0IrbHsm/VV++zk6et5ycLZmxXXgdue9pcDCyH3qlipXTQ/g3Dg3gduLNaae/AXi1nySeOmXQbW
f7YtKk26IBTZVjiT1kZXo/YJmheQrD6mdiOvqJwfKWlRamcmJTJw0wSv158p6RAiP2ftHJp9tG1w
VFeKtDU0m8RmhxU6FB6gpi9MGh76ZPdrlbI+pJ0+JQ6607980wlMEdM9iVe1vVmrqH+Qi70cxAwu
q2e6LY/RIysl8BeHCD7cK0uI6dW/C4ui3sSRv30v6C6y6iiZDtjIH8BnFnjsBXOZ0XRcQ9jmxTQC
ixa8LWkwDPfQ60KMkCtQ/OcUM0pDpD0gaO2GQjeDy9DNpgt40NjBN17Uup5r0GM2h5cEMqiXekr0
EJ95WJkDTrt+0e+RRCoAJDVUpZToHbVzPvYLU09qDR8M1ZJi3LNO3wHoxjimYI5qLzIu0WSwdqmd
lMi8Sy+ZcUE3tt51SuaCC41LasD8Q8295SfjF3P/ll7Yf5YykaiRPmES4QNBLiaLuYUfQOlBCpCq
AM+RBhtD9w8mmB3lhyTGHjlEYY8Hx05MV7V9h81A89q9K1vB1mnSqI2IoHBt8iyqY7tsHWSoNBbK
gL4xHMvL5XJ/40Ap7AXr5hKe0oAbzJ6mW5DPY/hImWJ9wmhiiqzxsM45VqrAKCh5+TuudhK3PBqY
2hA2pucobkYVdvXyv57tuwdzvdeUKvzA98PT/4cLjF5a/SFC2hhHIs1S0pGSNL7IFp0b+wPFaeW1
1lU11Xj5Cuyz8gbiMhT/Yh179j6f0u53CtROnVc+B3QHSX1ZSiymtmLnwTaNvnkXPbo+QVEk4936
+FJSJLvhpimIgETrXzYDZ8UnrL2064EZTdINm7LZ8H1HKUhmcw9AwAuxP1Kc1RubzJKI84Q2cJxI
/wJMKVJT1zVYqzfgTwbfIZ1z9WY/kFVG9KDcJPx+KoklocvSqCjnkWvvMvx95GQ7H80U+93dRUNv
LSr8i8nX5IZrtpA2HQHm1AwlArSUQe61vG+N1f0PLMQdQkm/+j2rb4DglSd5ElMRgTFDVwFjTnVH
J+llgalTr7dj8fYDQHBjkRZ+SVhyt0zofZzvQ1NuBWZgmShKOtJs/YIreVF692SDBWxRiPn7FgxD
8mT2XTycisU7tTk47CePzSJPimQb/k4g8u4cfvSkZjZ6nNqMJv/61RE/gATX2YuXo45RAHrJjTr6
6qDoePHG/4+0MJE8iEehT2eJji/kXzrXIpwR9cxdGDC8x/IREAvk6Kicz+dKzvsGT/Io/8eP0+Yg
14o14dBBEmytmyMYYnKs5loFG81gnPjz0qUEfAh1oXySQo8XUVAFctZ8U+q8MRaXBPqdXbjQ9P0H
qGiset/CWNa4IjM1sep7DE9ihD5J5Qhknt+lWCu0/kbXe5z9HSng/afB6+B46u+Cf4tHGCgFB3oS
YvrHMV5Qu2eVyyr/KHZvr4xFk23a0MPLvaFlT3qjiolBfxvip8ncIrA9TVk21L+kHggKt2K7Jaav
TQbHLYjhrl4expWQ82BILXWyqo4Y/NeiNcAUho3KdxTH1wEVa5DIu980/MmttPU7xIand3JKJa1H
L3Q/AjbYa0UI89QUWymZGus8JLHY8VWuTDq5ENiwbVzDhjSGkoaX2/cshi7P8Lk+/0FUV2q00cWT
gxa5r8UuDjbh6ucz1Hi5fTqpLqUC8lp/idHolHC7L1HwHVh+xjXzBU/Ek318DR9VbMBIeQTfUY0j
+NMydP6Kf9L2c0bGS+eisvuklSiqo7EyfYWJGKMWeo7GkCO4M5aXo41XqDqRhuCOkCtVMB+0Ya5o
012txFUIheyOFIYE1rv0mjly/QvGP872nVaRlyiVcujAkO+iTStNOELxNgZzMLBmJzq8+A9kVvE1
kf0Gbes9jVjwjFmWuVgkCulFpGQTy2gsb7hhSc0w7/pwXunWG1p1PWIe0Cbs23w+3YalXHB6udQ1
KHi87oxsc7ycyFNPdRUFxXA/K77lxGPGpt0LSAZi2RW7OPTl4dYxLUXTA3nBbv0mWhf6kkKHzvuo
wiTUMnVFe0rnUHlMU6edBp9BvdgXdCFNlbvFEvgZHzW1SpZ/aFi0mIeQ13vxJ8/ow457SUgJhBGK
6XMHBjCsL6EqSfPln8WefWoFM/znP74cWa6SHEpyBmnUYGdFm2Nh8yPICC+p9jSsSRtgI1DjimSz
PIe8sU3606ygzIXmTXIXTF5VdHx89oDG/ij1D7J/qtEjnyIgH9y95d9wGFmvAi8Kot2iKun78lQu
B0Rwb52/FTy85hCyk0bBJcnexYgqmp9OcY0yFWaCQ6IhpwqC5iwMwH5fgzEUfsYvX9KUR+ev4GC7
HUINa3wP+GwqPmUjJHwZwlEQWCk2XD55CoyKlKutstKjg7ASjcRhX1NWKpA/37qZmLMfO1SSZnky
JNZ6b4NOnJBpEWd3rCDfC1KyBSyQ+gyb2c8KX3N1nS79V+wi19DK/yRaXgkTofUF3hPkEzO9cb3o
0sKRZILNMTcTPhCYOV8XpzJiYPPrnLqdVjxfu66wEnvTd9O8ZMyHQ6yRlyz75Kf7VkWtgzLr3/Sm
aa3dZintSR/Z1lInpdWetZjvemMTyf5njfqwrVZSvP/k4aOSbMJ7fKNBmn+vNKiAKe5DAJq0Vpn6
2oPf6pAIOHxOe35gemDjqskRrPy5mB5Vo/UPrsOZQJyQcoFZWn+8widk6pR+8sbcSpTzpOprrzjW
JEbvuJyqCdbnge1M0CRzUSjmCaGkKn7GZg0ggA2mX3JA4qdVr9ONWKk83HDJDZcwIWyd8oBPkepN
ibS1S9N0B6Bp16CTGDpLpMtjwkxmjdJ/+JUJL7zHO2ftl2A5KnOfEuSjB/qg8/dCcmA5fg80tiv+
D2Aqp0rI4UrekhqpOH/GKd8rKhgtjbwYoio/hym4BOaW5DBq18JRoPPEy3OMz7jiY8zKO7o5PqHO
PKjm5b9qYdPm0SMsPedhwJPXhx+RKDy1FRuPOBYY64z+0NO7tIKd/FxruHFpxBntbWMpiLubZzM2
VabGThay83wr1YPkNCveK/fR2kB4WcRKefKb07vKdHyCzLVz3KFdywZClyJteiIN2VTLGcTge0Ae
GryNwnUd1qpuYbFeW56mTsNnmqj1Co5jY0g0Qv1pY4aZGD/D+AwnIjct0BLPYcv4ddrBXGwiXL5p
2mBsfUzSc+zfO4QJSNlG7xkyv9vzeT1li81WNmu2zyJZFa7L8tfnldEORWvLv2f5iAPX6MsbW3aR
ay7zLqCn6HVOSG4PubPOvmUkPBOvAIhSE02f7lUIRKYMWekdZ4flYIKPmeJLW3s/hEjiirhth/Fk
Ior0qasBz6zYFkx6JjT1yPjU3nMI7r/17Z7urlU8sL/8HlVrlgT/AFowIuUhyv4dgx9fV0fje3lB
n2gA0ZUMftrJIpOvca4bDRV4Q1zXESYJqdoTr0yaFeFOK449KMtmEyH5lNZkVJn/evLQWZ0409b5
+lgf+7kYs+kFAj/APpWzSlRibCwmGhCneeYrW7iHasHXknGwZ5l8/UknYScFTWjHYtbfFQS7XZ7n
AP3W/wAl+AMQyyCt80R4nXEcfSgClWDP39HRxTQtLPdw6nGXiYjk2nakyvZnpOFFYNRntTeQ5eq0
k4cEz7edO42SG0dv/7i/VBbS/sAgIbeMhaq9Y1JYy5RUdCywSYgBTMpQzPXJpq6yJkUN8NKgRp2k
j1qUyQRk5FWwHOghrTzq7mJj3OT4Y0B8CBFMehzXux9m4dxRCdk1H6UkUXGkXkuMQn6hYVZs9R7t
oC4M+tMxPL+vNGvk7pYo95N2YsvwSyLZ9t1o+mTQe41/omB4lit994YCs59rMXl8/ZfBxHIxvdBz
L6trPraIzkegipMhgsbIhk5WBE/dOpwugIO8f7K7lF70hBDtVrZlCU+588tzN4QVaqmhnWOqYq55
WpqrtGQ7skjAGQjPwA30wWIqCih34c3csRNwjNU1vCPmoAvj781rk39ly9bDHBOJoVuXCSdI5z/s
+GQQmIaaol4wHST4q64YUAcpQ+tCDGMpqZObEBx51TakGnHmqmrGOM7ivRYQB7bgcCKNGErfMYo7
sEfeFEqAPLraC4dNI+eITXOLRrcs8bbd5ehDFdTzErxxUVXagPsRXB1nFz8sCTfGBV3jlwszP0Y2
019kR1puHHy0YW1r7TuHezQxkc9HqLiiAIwDJp2iC3CxaVSey3Og1zV4wfxvaAfk4Fj0spi+kXK0
s95CXO9Hsja8zTQaIrcbCOV1LmcAGlTeC48GUWUETcyVl4yFct/tXzPmRBeIIcdPytMjUb36RavD
GziPehymrqzo71/k9dPVQ9IbSZzOiLKG4YbqmYx44VNrN4StwceXjnpvSv7jhGr88r1pafWGm972
XVnKcRN06z1nB3UJ3L3rrb/n7bQKTupZ36MqKgIK9r2yISZsKcXA/TSfIIWUaEyHWYsl3DMGEta0
zdtXbAw3/d5YuYAn1MdIObdNGqkIQoHDSgyb5ETh2to+WwhicUY0XRQsg+xqsf0ScL4D0gkQiJGG
8kRyuQUhoPwKs1FSRaQedFlPGgoOIwixsyzETco1WO+4Hp4qM8gWQ3eNLDlYZJXHdcrdpTLylafH
59J+bbTnS7bc31n3Ty+L4o5cHBZSpUCqPUg+mEt4kro2pY2ZrCQKL1/jhYTpPf5gQofHRGfUEAdD
x81hlPEAXFzZxS/cyJGQnvdB4OIr63pmplSJTnXCE+mX2YZcdgaS+ujY7trYo796enLZ9wJeJIY/
AF6287E4WVK5zTdD06zEVkxWVYOM+ZpzKj1YGn97nMCrIh0VC/IYgfzvcVQ1au7t1XHx3pWvpbRx
Y/+YiRdiJHUeso02CkhIkBdpOB1FPiNzKOOU8raOPRN5+yKLbKHD9WOHfAqosAQVzsKeADqBU/6a
GYl2OI3RFKF7URuPg614MNP6irObOMW9KwDDhtush2rUW9QliNWyqhOXJsreQVZBYikaXDL8K8AO
RqtthfuU/OQnkhUtVQ5dyvyFhRqdzZ4viDCmsnQs9ROBNfouKSJxCc1JyCroSzYU7fMLSAmN9WIe
tSgSD6aaqFprRTRjZ08yjaCQRLtaVvZSr3UATJcdzJAzuqQeFXCn/wooup5wuf4JnXzy58HOcXkb
I05E1I2zprX8kr9J3ZgM6kDwqpCmQqQBXmuvLLkSP9bzwBAB2OemtOTqr6lcfHimW5xxx1TjibZo
AMlDdse+ppWVw2amuu5zXs4bsdB/mOXNHVwFJW8AYle/8sGBBli/XVKY5WfZR1uewbUhjXhy/yyD
ub5orP0e98e6Q61l5FaSloQBWaVLUtWyFd3hEVbP/M06El1wGjD7Ze0cdNzShfxwFKG5BkTq3QC8
paSzpMCbeVjY4UMoXmrIbPtIJ0ON/F0gyKRw9LI6UmeU32xzUpcVEd/VzHpMYR0eii3+fJ4J8U5C
GQvjzi5u1nzpYExfdoQLBZFQK4nBBig3QOALpq1luvDfUm0SjpFuHN3JcdOLOqj2Qg1PXToFhcKY
jZvWri3NKlxlQ/1kyE/WXNdUqDOvFiBDbFPall52KVn9z8WMSVNkSbWvfupB0FHvbmuFpi+7usP2
Rg1Nin9KTR2rwq0SPjlAQDKvSkgJg3S1Yev+JdPZ9nSyudFnmseNhiSKeuFmGhpnPWKIaFaZFpoh
R4EUPAObC7QGQtUkKEQCJbGin3+ZdMgn1rLQBrSOXkMJkoce00TYfMA7dUP99jESlzph8owb3vs1
ZSo7uCJ+q30AF+TXJ1lpLV3Slgxl8eWN8xgQF3deJ2gmZQpsFuM/AFRUpN/MhZKVNpHQAdq3nCDW
q7AKwLDPohOHX+vVX7gn80M1IlVysslkFT3MuTCVWaOe+67AWCYr7fGfY4IlPaQ9Q9vAuKnrpMbt
7Jefd4u3bPg1ey0BFn7J0dciXGyuDh09g5GdLBHYvNpvaM3Ee1+FxeRcULb/QUAedytV9KtmNhQt
Ef4gWNlpSiUdTS6u1eli6D2C5wtPmjXYqMn2UT1iD7Xj0z01uusap4LlKhg17rqheit69bLq56js
LM2xHqaXeGtnQjHYPOFeq3eWRFjl9kgMdVL+CZV+q69IeuPjVv2gN/cxyhZ0BeQLrCuipdGTOaDm
ZQkVFX/n2UgTaBwwnB8oymw5ywTWzyWq0B+/7jcoekUU4Vq3GQG+oZGdf5mvBRG1gSXVL3okG1WK
bIzzG3GyFS88NCoSmdFxYCGFIVUclGO250w8ILaPPPgtURvLpaxZxMZ+54HyWh+XsQPopHQNVBjX
j0tCBv5OuFAIy2rr+aYNVWhG1wgHS4T18+VpHQSbR5FWx4WJjjNunoU2kRbUH0uz4kMSlvriXWPq
v2uiZTdNMHL7eXUp9gN13ZpY5q0SpzpOcFCLraJAl93EkiwiPQ8GpemamtpzZ10NCSBC689pUBIq
S9ybbfAWMudmjV/QxQHt5j1yJDMkpotngjRzYMvbP2XAMAlyCU+KLuQZMXoAkfbNYwsO1/J4dSX9
hIuyIMsGt76UT/K5AQtHbPAZiO8wpitsTN0UFDv43/YdySosFrUmriqoHdANGkGf/ZUhWQ1LJF4O
dG0CVXiovJ/SeuoXH2lpZV7qzpcSq7iUwKN5kkqTtlBqQJOJ+OxRVIqJrINPYXN1iCeaG2KDSoU+
2knwuCYDig0QXmok2hIFiTTlFy+zE9oExVNbYnbmM9Ga8Pcp0sfvhFHDT5YJhCbPAS4PxdKr1n/T
2VDLdiALbetNhr51k6QATLWzYxjUX9xJee1ORlUOjvF9nXdIBCb6i15oDhUT7oLdSTMhdvbfvSLe
UfF10i6HOtqGJdjHSasRI7HplkoQigJOGWBAgqMxfuyOigejKwaaKwv2lnyPAwbBgTBEuftDIMaR
VT/RVUJXewsGoheg+yg0StcjK1SCsIfAnMCULA5CPUSbyEeRk57yCmk+Sr1y6GUEfOW/z785Mz41
wocDKR37vqZkJOew64Kkyql6sfSSXW3HRogRgdx63AH9kAqwSBeosO08RDGQ14P9E7KhzutBzcaa
uv1uAykHz/P9or360YimpVXwWiLxmOABohREbOlQlkiMQub98YFYVR952nV1mRsWVGNCQ3dj5iVr
pUs0gU1GtuXRJ8TVsBRiWQ+GoiNAuepq5iAMLSBfSZket30F25KgopnROkGPAdFKd9v3GAdNFYqE
1TsWSYgut90Ao+Y6AmfAEZfGEb7n1xm9ftwb5MKU/QZadRfNwPvu4B7vcAYQx2VS0LybQ933tXTv
0cercMbZWdYYRZM0Ef6myP/bSZ9I6E/71AspA6+VCczOIAgEUc2Q+JEnBBg4dc/nU61c7nf76IkV
6AArXuPmj9nGH+1yo7OlyUHiVHg72I4yQU6katuFR67MwkUkPAZVAh/alsingK6LKztbYVoHV3W4
3eVs278UquzjFWgYuZqUt55WNx2uoEzyMMkvEM84kND8Xvw6PL8j6k0TtndX66cpDYRkZRW0leTS
E0aHq52Po5yvIFE1QdvXTDDgITeHVbGI+mm2mte/2jF80mVO8y945lhJkOhyfMKbOOVRv4LV23Zj
PNfHnIdC/5LedBCQSvlIIvOIfWv8Mv706SafFEoIxO5LCO3G26IWzoq+Npr8/TSMc13GYGJHNUnC
yWGGdx2jJtmltYcQPKrBGqh2dKSf2SyMPdGWLBLJ7uY2k1xKFnwhrE4SeLMQ90t/a06akHlSyQo/
0XTGiQzq6OgELS6DuT/dNwGCOmDGaqp9CRuTmTF5H7TsEXGahzt7nKXDlra1fP5REIcW0KVgTypl
vyfszIoD474TcXYhngLx3xXyVEuCAIhGRsr8nohMno/8tKZHE81skY1WoyIPqu6KugIKA4Wg72g9
Kc1INIrno83lxQiFo9sxLGuRrnuk491p4jHZY0Mjipam/fzL9FAQxkUSdfCBW+jN937KyHCs+T4f
+cBgWyK5ZRouloP3jOS0+lEbSaEEtAUmlWb4Kkhn8oT310yxvDIVv2W1MY89rZLb9O5/ct6ubwVA
MYO0yp+1rQPr6nx+2FUuNyMsfqaFc55Zojnjfp5N4YfNDxjSHKBboGBLpLwj4Fu4Z1RfAJuHEoxY
2yrojm0m0SyONBj7Uc2zDfTzT6oJDiw+eMGterzBwspzpYpAR6Vn0ApI1iArnmCfwuZ11x5OSmo5
Fw0o0jGLojgD4zMOP8Yvd422TPbYl1FaFxRFUNR7JHonGWc20cVHCqANg1vgeThREs9HVTCznNA7
K6rG4odsD9EI16Fdak4P2oLfcISVNjsetF97eHx1XdFgTV8+2tGpe8szRdVzaD7SLMr+5Curj/R/
wIXSRK+1stm4y07dAaQdwy97kkX0MQx7+lZxCBvko3T32hQt/EY8tmCxRhaaKwVhOtHxge7v/n82
xqGrVujY1Xp+QpPSbmvaYEn5oGh/xQiikxg9zEk16kD+AvxX+jy/jvc0tR11aGvdP9k1EeGbF4/e
rNSalgEQyMjARcvreSKlJjbbyV9VrzNeztIh6AviXMP38PurU+MhmDP520Tizz2O/q0fLmlqpN+8
s89fuTp52ebzm4l1pNuGdsiY4keOEeuyd3ZsVLE7Pk99FZcvh+n/6dosv6qvpD4wPWgRQhvN45Sf
VYYgLoyO8N2ebiVCvGcSQkkGhKI1ADcNOu2sA8Wk8+gm5z5YozWzYon4ryqRR3WvJbC5gSjAK6+A
MmgicBsCiIi5eGWWnf1F1Buv2cZSq1CQiATSgf0NRape499LPIv0/SMfAGSRoy9C9xGCoqlNtXCJ
nUiF4FwyvKJrg4usZ4JTsnS4dD/btUhZa3H+IuS1iMPZV7JregNxxS/tlB/M9GPwbgOOpNHwB49D
wU3tMOa1boscUTOT9FtT1NBMPuPRc/HVoAEChRyVRukbwbaLuWkUw5vNIL8UVP+bzxrVZL9WhfOo
OuzWFQkIYXr09gBskGkhCmtjYJ6bdl5VWU1yn86PJu4cLgFdH3XJ3N8KebkW/uOms/RU7+A0kPnu
oTyUe+5/UJOgZpnKmxzkgCbPt25lhFYIey2rXwDi9cx8eK8twv/B4SZXvd7otmJK+GlQQ/3blrVt
p7YYWEsEyvI8+wdwKEspQTKzbzxB36BV8NSZM3Jssdui96EXBK7yrjLb1XEpY+pE6wMA1tOi0PD7
ZS8NZmYVxHocMeZEnoie573NiboXo+oZj/M7TfTSIVeMsbqq0YydTkPDLwPZFnKknNONTf5uKhE2
59QiyIBL2uIEq1sCmHA7xAgSl1RHD9+c3gyxEDxci/3RMZGLaq2RyxRhUjsfev5LRGEA8nxiRpch
iF61KcLp3CmQGunAqv50h1bjF7swrGu7rYWQ31NtiE9NaFGIJ0NPemMuUsQM6GSK227HTi/JpN4K
MTdljKvQRWWgBTx3wEMNx3V3PhR8YrXLOgm+aFkuY7WWIcVKdmVjqShyuUErEqa6xXKAjwbalaeq
XuUwBemo5OZ58KroDp70N++/0XIkTOkpwbJ/WOkbxZmLXIYO3psKQI2lUKDnQQ/3azEfbUnnZjF4
JGIE0Vo+gSwPmEswYYduJ2VdqxN7g8s8eL2LH5w8d/4UeqnzaI948OUE7XEn0D1+yuh8KkaNbGhC
hZY+PYrwsecDrIEWKmFfnwFG1iY+0eHgcXg2jVrwUHMDKaf1+Q/uUwwnHt4HBMbi+exJqhYOTb6h
4Ha7hSHn0SKzwyAC8ZWaaThP3KI6spywpPYeGwc33n+0chY2AgvgoenoKES+q6IIyG9dn6sCtQl8
gngLeWILp8euBKI/OYJn6RH9vnVDVM2CZgs751OnQrErTypVQMcI9aYkJ5sg4Nnrqcm3hIrDJjst
mLnQIaeItEufJZq28cwclN64/vYeT0TMX4xQhBKixWtbHqNTe8/HXZtjpL3ig20wM5u9EjDxphvu
PYHJZJGEVAC0HTWWJm76Ci/hn8QrU971tvH5hmBy1vkIesFWaa7xMvkfAd+PNEuNeefawueYkBCN
1j7VUF0MeH8NeUA+FmNHkjHlSfOxg8uAzlLPhKlXuEOqD0TApbo/Y14YDwxHVo4LPkbr9eS3CEtD
Yb4Pz02nE0OwoKXWJpWonjnPwPkD3xT8FlDX8naAomOFqJ0aWs4TJNSjLOeQmTjjQNJwccfxk24G
YO3R+glAVzdtheMkYfehR6ZoWuIczHkxDWgsi+hx2FYMS+ygwNJG6CIAQnhPaBbfk7cec5v71KQq
QF8TzQPYTpm9ZLrG+b3KfRLHOwcbKQ2dSgXKjVAl8K4fHm7+sIlirxDhd1Ms2P8sA5aa9Qt5GZ9p
h8MbDay8opjnvhGEGJQFtj95NV8lAH2u9FhlHvhK/kdexh/Afd1lOzif1s38nwwHIQ3nl/zXkHtE
whWbOvDf+Yt1gq33FetUu6dxIz6GMcvpc/J0voNPjc21TuGLW82TjUQJ/D5LNUYmfIorSuyHP8pW
HOLPryXQQkSjF097r/X1cN+ApV0Y62Zgm1aZwmLYdBE9IBHMig+XMdiisUIACISZZL673LOLJd0b
PzGdLF76s990VtoYfH21gTWosaoy13ZblEAjAu/x77D4jZrnBySnh5V0f9irqA3h6OLmLlixydK2
Km8V0/eLQJCJd2UunnQuFH1FW6SV4FVZVgK45oKTeb2vtxFEsOAT1BepKHnPqY8YKQpXyYVGYuDb
lJx2qTc3UoGoRepy/dQjgBiqTohBp9vGsBC4iDoqgIRB6SHuS7pBUQbolmA2eYK+1RbizuMhfZD1
Yimw3J0wNecWkCznvagw6f++utOG+jN6+D8aSlD+7PM/0H14387Cdgotx6YuEzMYkWfjLPaXnugu
7WGhsz5DwdBoq2LppWE3pFfGWsL7mcrXLxBjUZ7svHkMQQHWdn/wEaKaPZ0Kfl9WgR1MSNuaAYyn
veJIXOEQyUXHn2ktGkDjVc0ZJMZP+MjGJTrBCIX5HPN5ORzARfle4PRMI3/cEMrinEL7pPrQcgAm
QRcG5sRm9nzvz7LTGd35EsXn1jO+ZbqSsIMUfniDbiLWo43LAaqUImu4GMBu+D9MZBI4p7GxGBPU
9qXJgd510lDMqkBdsRTufEzuh6KxIEtEHc+MB4cusUSyjdvWEItc2b52dk1PJ09BCS4xgJm95yV2
oLA05c7ydY9IN7c0uqDC3WXUoZOVMSAzFOynqfYS/JhXRpjXDY2cxHQW1lWY3iEMOI5z2K4E40Am
bxkgRBvjkknupL8E3v1nHphZDw21iznI4lrtFsBVMCWFnks78sG+8/pbbzu8LJ2cxfsZ9TrPUCCJ
fNOrildR9K2GZhl4e2ItlcdI77uybcK0ctYV/z32LyqFRwkUF370mOaNTJDnApQKD+cd7Hh8Vt6s
BgjtiXhyJxFC4mDLbheTTJADCgH/EK2nFNFxastcHxuebTG1CmvfZiHHZZuAmt6mBA7ud45egAEH
6vSeRA690cK6VKwYryJMTCMzXeU6XrgDcZd647LaL29+igBUvw5AJAcCMXOdB7z1H5qPfr7aHoCX
a0ZGYYOcgwhnJ2kxmcVxiIckr6we9SMisrLDNja9vPrL3evH8yovV12hCxQO2CMX3jRsbfuYs+vn
x4fmDGRue+aU5sxbR7oNvhZUBngvlDnq1z2coN3uXaTcqHDuQ8FSwO2JQPtlVWbTjXZUXvqllvUG
zs0YkpjkA4nzb25F/hBD3DFwrdyWlNzvIpKPnI9VQxvLNSJ1fqu8dR8dzKSYqBd3I5V/+ZqZaL6p
XORxas6noT6ocF04dmbfIU1T8c3U+5wRm20A6VfniHfPL6QjKvc17thf5+EocjygnPWWpXgfXEFN
42mQb+sr/F/tBvWHPodBn6sv8tEyjja1AA8Cbf8nGdWyoJf5PXBBo1jjFNyAZO1QrSab9x0TamC2
ehEgh0zZxzztTg36oRXpvr0ihnFX5213cTbXQY/N7MK3K/c4E9Jlqmvw8O1wIgPAQi7MsZebwN7E
HnuCiT3WDQTftZCIVk98UXsniAt2r1ph6hqad5V/LwA6DqkS5dA+wdGF8LXDrEQI4bmiojxxkxHn
XNlXpBvU2zrC22zC5T+eHEgatzqie3LSm/2nRp2hFhItciBU6T97+frOJIznl5bEEUDI9WfusIad
rk2Q8ak4Ean+B3vetX83RUiFqT4/R3D68AKcf2FLgg8A3KOOxNI9ioClXsMRhP1Az9s2UKUCk+Kz
LcS/XDKNTjAwDwVlVnhoUX9EnCeRr5YlXJ+g9/To1V3IndEhcP2yGcjAYxPxySIQIy0m5EDVge1l
kitc7uh9GXU0KRiJqtLP5VUT3qUJxpKYRSkH7WyXH2m1L3yyLkEFgUbObR5Jq9x3AUGa9kA6jb6P
KTWbHC3u73dglGko901Xx4ksSPFL83ue9DDiofjEZ/NmHiIrr5J/8kFqolNOv4jiGyUwtgMicwSN
N5OFFRM+yuBA1yy19rn+p271qFonVuXoz9ZhhtQuKf/paf98LNeZB2wWsSM+OhdZdYjCUgT73XS5
t4vJBv+/WnkzSZUl+2F+AMtlgGrlp94+lo9/qE8XTyiFpFV9gbOD6jMcN7vzcjGvj2VT3IK+hPtj
T8qrAEMcBUNamFAGySP2ooPl1alf/JInO12y3/s9xDVROvNKoPPOHW1lbf+pJpKXf3HS5S7da9vy
INWAwYUPp1urFTYS85+n2fmxx1xFPfGBVhea74L+AK0SuyP9oqj3tOiAenXsgWrKxNx/dLafNUo5
+YTCGGRK9sq6Hg+OG8sA/a8BTBtK/CIp6PFAcNy1VkHa5XWRd5vjzYli1npq6wL7sAkUWVVNpPPJ
vEfQzyxMG5DdjoC7s8mNMorWbTvIFeizUvxZnp9clWIpMp69WpnlIIxSDKL7JZ5VV7Uydg9sMClI
6OuJJOrHBMGEd9LJFJhMEMPTsVrDc/RzzXTX4mmsMsOgueOSnWx6xb1kaqNckiRCEkBlsgYQXwm8
IgMdREXmrGEknJ1vxSFgKpjvXJPRHNKLg4vF2igMCsC8KYB2ZlIpro3t1p3oFI17MD9ljuLttJhv
VqyyfOl6xTXB+nAfFsgW4nDmzsxZ+acCsUb+bov4QWytpNqqeB0STBNYCZnqy+PhvHaG4PUaNDMO
aXSth5qqLXOAiqdhX/+Bc6ivrfNVq/B0hfLOGaAu4wg3wLMq0+yY9LznPfWEflXDXtxCT/GRDtiv
Lbx03/F/7d0J9vglzAJmYsnWUx0UMHCoCEiizASTWN2UPtWFdmTlYKrQEMbbROcj+8JdYRdNTPSI
cmilsE4kIboqH0Q8VKFppxhBOkK/asdk4oXFSiVijBtwp5KCi2D82Uq9WW1nthwSVp7NLmN2C8JY
vFoEkkmea0D95VhZKdpQnFA9l4RzCjeg/JSKFNmORQc5G0/j/4371LHCc81XSYWdFRH9IaT+KVz/
jAz+eIzrZFERQNc6WtvvwPYmBswBAfkdGMTEV0N5gHCUOKRFB5MpuE+t1N1G3ut9lFMm2tGISPn+
t2ROKksAfOZmntpALCeWiO7HW1dpioQ4q2oK5I2YtH/dNUrCC2kKPIfdUwkCex8F2l/SzDDdtG78
QQJIW3avNLxmda1kEyQsxyW7hOSWnCvobx/J5WkaTp5eBorpLWHuuZeEabcQO9boOQu7cfl5ViiO
tfjl9PfIqpU40ibcEV6spwTEZ03bh8UgbIgikAkXz6jgG7gw4DKov4ft2/YMRDoBnGJOwwhw76o/
fXLncw8RE9OfGB28Yh8zJ62BsVvnKfAZGR7JX3sL6YzrfJ82OdHPSBkHg0doO+EiDbd+ejVQxptn
9/hyouoQhp0M7VXnNH3xHdh7A/XfsMN73KpM5c8kl6lWBVPpZxy8nDo48diTw67u4t883Hqa0Sla
wKH4bH9InSmVKS+ML1ycrPriFin55Wbk9WHjhsZvUyhHBG6g6DjX4ekLlz3JzitidkXx6tt1KkyD
oiKlUJsaiZ8TV759fShoCjDGDoTCdtJ2F53piLGiJy2tuA4WB6rZMemPWq/p9NUN5/uQmfNO0t9k
R2VOqRwr+l/9hN3moa5RFI/Ln+6k0KgWo1ctpstNgIPgAVMmFrzVA3upFsxKhu110b8C6ILHXobp
rziNKV6qUcG+VZwzx8/Ew4Dg6Uhy2I8YUuwbkSI/tCx4utfotrN39WscLVmfxLS/yR4xGOyURh3X
zPDc0Sk8PAf9JQY9cgKAhl6Xbb3eoHULZwbrE0xLdUPahpWaKvjRrt1StNYjDDHA1cbCjNwevSgP
T/ROdQaK589SLWBySq6lVzKec328RhFwVTJQZEGL58DCXeTmbmzEpoE//pjRDRw/nIatpFrYxJx6
/q7f3w+0M9iTxMfBzxz9T+b635G9AqPYiSrdxPZa5fKJCDBT5JLIsoHRM1aUL8hJu18jkbOX9JEj
69tnHptwCHY2o73b5D76M1MUox8AYOKBWEPV81nV1+HWCikcKtdobfR8ku+38qXPrkOB6s5panFC
zuDJ5kdgxpAsBnjDvhT+a/biusGyH4P2dEaoj97auGoWA/tGhRLtnfbdqJI1o2QMAV1zUowvMJ1c
CYci5Mu0Hw78B/5eVdB2rQrEjtmRWddC5WjI8Ps3kTDV6kh0QIJFo0drX/FzQWPjhCECJjZCs75a
Y1jWLOtxlRDaTDv083SdbK20OjRUgFnfnVHbO8TK9/lWqaZY9ub45XkCHIehMDs9W/dfFmFUWK37
0uV1xi4GNKjDlXsyf94NKhONfyUPJhx9uk+33U+zNE/rHbu3N7cbF7gLEBT/H9rtEkJSzFQWc30P
+phSgNQ++QUEXmWE90sKM2pkCMkf13U8LoIw85i5RIKq2hYEpDrE0CM6bQYAZjuRttt7L6IPr+jO
7S2qnnU7bG7PIVThBs6I5A5cALu4+YxQ6mYOzwninbocySMPW/twUY/q1rM8GVXTMym9n0DTK7U9
XP/GOEU++/0F974Fr1K7dusTkOY79ItsUoSeXxqKqrIRpsSdk19urP2ePeERVcOB/xdanDLbFXaN
BPzUpDJ6HqC9t3qNX6Z8Hi2X3OSp42YUN0Tnoo0c+gpOnbdAt2WGyfWSGJo9JAPR6kphswkGA+06
izjLlXfPqKahpDNtrvdg8gL1Wd81dSvbCSkF+K6398oh3tHxklIdW7ClXvbMBvoyWPCGzKlZna5z
/oodnXa+Bc1XprqMgT3U1wGWeKHysI/9PMTVH8OqwCU5zwe1/DU8GEMbcRyYiZxjF2gwAWQGkFk8
E8XYaZi9ReaNfd2utXX+nkopTvBgN2kcHXK2yFrXHmroJSRaJdzfj+bJ4ey8bG7JFU+d7cAJJoCk
8/CHyt8a3NpecdGT6kvJswQdxaQ7YnjRSj/M/yvfbFWpIFsl7ZM8FSD3siOz7SArxNf4I5r07Lh4
shuyCbTWimvokPeZNhc6SYTYGkdKwtJVvWAcnF8AGzGF8ww4c7lHX8rXnjwDEod+dtQtBlbO80Hq
QPdzSh3b0tW3Y6sMaQjvApVLPq0fE6hGGSjK12kmhCVWb2CqSklaNXhvMYTx8g5HPGjgelzOf7xq
PFSmEpcWqud3+sbCO/cL9QSYQadcDdWm75IymU956ooSqpSchMOvsSkRdmmjBhttanyxOWFsH1H9
mB3jGBXwNemv7A4HpAotJ1vCBkscks1s6RbTz/nZSmFj29SIAHK95RB25nPxwQyKH7g9Th550g+k
FExn6y1Os680k+MMQM3id82zXJ/ibO6uFID0VxleMRImUptOzsU6oGTnp+67FSTbEMpMK04UDA0E
cW25ryBVMKo0mngWkChHcjiqErj00whGoA8RavBtqKJz3bQl1cNuUHfvD1s3cCMQnmaTY5PSlDEE
ElkDSaZMozqKCI+LAJPO8aSMLIT6j6SpfJnOLphK0E/S849vWpZZj3uJ5/XQMmlVcKUH/xOdt9o+
cSw32JkWdjmO7GhC2GH7tIrZaynxq8DWi8jbBVzwOFAKNpGsENt1kNcrdnDKVZ91eviw6drEfOox
8enBv6S49tAekkJx+hgjnCbmvF+cAXuQDmuOTkLBztM1GZIBfATgz5pnrD/vFhnGUmN33fQmOz9y
XbDyzXYxhmemDz9FSgTRaGJIu/irxqzOfej4ob2grlAHxzs6Ri/m706afmzhnuXx2F04kx4XVoI7
7rkajGW4Jeoju9qQIaOEQJUbbHRaVB4ETIVOelFSbHIE1Rk6rSa/FRiXsPKfXvJ6jWGKJtQSYcPv
I/sK1pGWlMwF49mkLrKNQA38KL0rJMwlmQ8FL+FDEmX2UjyV0FO7M2OBoiD+xS8guvKpvhvIutKL
16fbhIBdbQJvnSvVaSv1wkF6U17ul3NoapEt2lL+dHZ+/hwg2AOxYmhswH3XZcISHW0vAfQLvHjM
7K6L+uimzqgv+a4rBH+YlVGkbHqejs9t/citA0/63+KCcA+22gE+ukWlApY68/3HyboVuYDTMGm+
hQlFuqvpmc9Cwr1IttGYCdpAHErx7imMryE6YR/BvkqbVaprSMpY2O0odwnwq2b+vHcGajlO1uVH
y+iCSY+GYV/EN7n/PXG3s4ZohX4qHAawyeTOHzmMKVS2R92l12OQOjeX7rArI/dY1KZDQTiQGUXn
ZIO0Ek66plDz8iwRNgmL1cCSUM+G1Tg8Gr4irQ7/aAj8o/QddKlmH/RvtCUigp+aUD8EdszlASJu
3BIbRms52FTMbkWX7Sot+3WQvnA2AGM2FU1qdmou9W9FvSREl/khFxqK1WmaLm1P3rORJy9u99lq
XV63MrsJGishlNLwelY716Z3V21Hn6wUmIl2zSYfjOPKpXiWS2DII+yC3IjhqBkBRPIDuV3rcSQp
03xuoJnqB2+lT6NU3mionK0iEb1pdam+/sXp45mE0lTbewLQBmIrc+KJu6Euqsb2nSNPN/p6WROp
QruiCC7+ltLQJ5b5hxxL9D1h12rLr6KlyB+UxwQTRa8Wjmifs0qNUBaNsyLU6DPsY2P/AliT/PTd
Y8sbP3ff6W0wVguM+6/x4kkVOTG9ujW8EjPDSDMPKaVMKi5AQgsNCsH+e4VJ+kXWB8leDb93tgQP
xP4nkIh333iivISxCeq08T1xwKhe/fLp0MXCLPVt78qqr6UBOtflzq9rnpXsVQT5179vyjUpu06Z
5xpc9+6rHcX4NlTa1OPJAKr6G37Hl9E6Ddkg7XlGIqjPnCcJ5T6SBNmmrb8jzIAvOqz8XrVpcgVc
N/CeJpKcz0C7PEr6OCYs/ZHQj1bTyDyKXrUSfygb4TFwvFj66VBEJ2fpqSNjhRiOvycuFynL64FE
N24vb2J8D8GKJJyFHeg2jEHNN1wSdVxHzr6m0ol5c6VCogQtmaSKrv5pq9m/lZ38YVgA56KxkhHx
bSWNuwpDFxy9UM4hdWq0ZP1Jrn0Da3AWr2hp5jKrNNzjKfAPM+xX9n9cp/epaAvHYXjvgggov2vp
mocKLTMBbFss0XGA9TcY/AeP62++RZkaQkIDpNkWVlJUdP26K7iWslwzl0T/A18OsecmCUYGsiVH
mjBOINzx6hoUDSglY0sKNT9Mjg823nY159tSnG03BWqPRoxHjrtQKnpYsmZH8tX2OHyj1Cfe+c8W
0nACi59/MRJ90YU7lnRGBaZWXGu7PNRPKeDoCThyspuETZhlfaWwX33Fd8Nf2pkMBV34MrWtMWZH
2I7na6e3b7X0WSM7RprW35UIXvedTvOF2RWWPuD8BOLj7FHX+qNa/Y1L2nZGcr8VNt8BTT/SSZ2u
ZInZRScDJf25HbKFgmtjT5X1cEP3N0kr2NymPXq5LpqhJUdfjhrWqr/ezZb9Uq/Yt76gFALgPsK1
c+b/lST4WQgVyRgk6SRBh1XiCTfMg0GaF85rESMdJpRQuVkzm5BfaubCzWa4uOfZazxTI8xv21t2
2SIdTQhK0gxTd/VnxYo0vJmt2mTalfoAtQpqt1cs0XA+aFuIs+5uipRR2Hv+kxKjXhbto0mp9ASL
LPXGI9B2b1csvWW0eDh/shJNDcSU458l8WgLslNoRO/p1JpM3AMnHG/XDahX9BXVrNmQTu3CJfIZ
bVx5j2ENLrJFKl7a4X/HfZingEPappcfaHvbzjByb5RnC/v2ZYt+Ekrv8QwHxccfoetL8qGr2cyK
B9ac5Wh0/iBQEBU7wZaN742AJ1vy4xmhCl+4WKZHlavItuczWxcLOnQee+/CpFk9J9bXAJ3EJ6Ly
+PJgdnNGNdOjxydMtDH4ILO/r0Y5+xa5ogKefG3knyiM7S0L9WYdhEo1ynSA9PR3x8wuHFlNvlSI
QpU/U6BHXpZYH/IubdC+cm6VUVyYTZg2dQomrIjgatE0PmyshByZ8OBv4oXrCZ2c1SUOYPgU+GC7
uSGXZo6qTp03BNaEXrTwnxHr63bCoA6XNbtBSoiM5AEjCCwttxu/IsdTy0j5PCIHebS20LWhm88k
WZgMXZSW/m6hAz5dDb7AG6dHoE5dIU38JKHE5S1OFw3Pnu+OnUOl8Y7sRnpFeXAXJg9bXwjhhTjO
Gz6JjGE0kdbiCeoVGTMkj1uhp8KxTBgvSTWtbrLZY2wbr+X/wMHdMppr083tUL4btgD12bVwko2l
yqbI3lQdsVJ2ULr/0pIRksa0tSL3lK/Dc5pDeiuk7QDYoNfEeUmZPiS+1jeUSlXmzGBwqGpooT80
IsQ1pXjiBNX8TqzgDakRE51XFykxAi2vhkTg1x0dXwAPclQ0MqyldqhpKq0vLqbYv1/sKFz0dugb
0yz9G3CpS1gwx+OhwVV6djRrJSGUGAcFIOzGOx189dBtkg7Ojq98WWaryqvCG9NdwvVLZYeqLgLE
4YaUWj/cLuB5qEcmDIaRl4STCWwEEVKEAMQjRvF8gIKUbk2gH0umv2qAC9jOra9l1ALP7GgcSb1z
4IYL4matsBw4QFth2wbdfZp7gVkW3o+iXfeCzWybr7vj6yqDhUfzL1CZ30KlEJzJNk17tdJOfYpS
NPSMn3haX00N9/wjiED0LIYYUANQxccuGeZLtLhU+SC58z/LPxQuVcFDQ50tEbPzsTzafajKf49a
N+EIpqFBf3iIB7kWXUe7hbT8Qwpu33WT4UAuIECst+lzSvjIserWpXPMTEBjH+qQbSamSElJD6uz
1bRQ6/lBTyAgoF3C78igqZfiDrXoUjJRbgeBgF5wXol7x2iDLIgGD8oszTqiNgn9d0YImpWLhSXm
sP1BgDap8J/wcrI5o+LPGx8EedagPVuNkN7wtUx5tsyRE2HnxGGfsGFmd5okQWJ8XXKognkUVTJz
qnvsjkWcHiuuoYQ0WlCKpYGyeyvahXDdnQV4jeNyFzxmq5dpQj1QqvT/KsY64Qavbzr+n2oSgLrY
wIuxt7Cjttg2FaSpA7ZcG82tcn3I8/z1eBGnfExGw3zJ3VCwF4OBq8o5TaS8Uhlw7571JYUREDb/
O8qY435RmEzC/81GEHQ75KeRZRVMY0ShYcuKSgV4n+0odk60KOKWel5p4FGnqYgM+zVb0HP07aPp
PABnk54jDSe+QB7tVpgf4JnV0OaYEzN7q+hkjsxFYFJCIu3Mt/oRupCihn/H9ky4LJPa0qpDzVJ5
nT205kwsi1FL78meBKcwliOWd+MaeWoAzcjR4QGkzPuYEBidF348k1wuvN65S/D7BnlBelKatL/Z
ZPfUV8cBOA6CaXcrVMCXN6AlMYe++jhm2OTLdqc/81rwMsYB4+7UVwOP+OYSOkuSw+hWuc6YlKbh
2QeCVshgVY6yumazZ+AMZSg7uCl1OL7NO7eA5Zc66e6WyenDS1t57r0fl3X0l1ml8bPxQ+mp3Y7I
tt3ut0RMbUOhDys/CvhSVQexRddLeM73drAmeuZCcDFmJPSqLUL8sdt15e2PS4DUuLMETB7f3KZN
oWOjSwXt7ilDPZl/dWpoS/pWTmsOvBUxAWiqEFSrEfONRhNxCvFcJBonAp2bKVmiim3pvGxiwn9h
HR4H1xs61JIiex2ySEOmVYc2ReXbMnd6lfPtYJUSnDhPnTud6VjBE7hXgHlNRN8FpV7As+aDBucf
Q/96z9EUlGOYEll7eS/1m1CSMQzu0rpN5Gxo6qNZOfaHBmN3t37zM7sYGfPnZHpHdWV705WzSW88
fMHfJJVXY+1QH46aPHrvWeR9+nIcoZLDNx5uP35evpBRNjzDz0WAn+bHT+XPoDqNo8cLopUznSrb
e8+mAMLJ6swA9C/Ddg7X7qVq7OcLgrj3btXf3/blQZOS+pmlEe0+muirS0MHsQs5xyx25StsqctV
ieY0ZwOONzNgvJHOP+dD+tbiNrYcx57h6Q/y5TKCYjvRCy2XAf19fg7NbZxyjcvGGvVUhf8OaI3o
ccJVjCqjrPorYQRuVCY8BaZ+iiEBpddcGn6dJpCsg4zfd/Vw8ybiZlgsZqqBiN3sXi9NxQqU2Pmr
Z5e9f24hiQjGyYbQ0KyyTehEK/aKTPhm0p2r/U7IpnyFbiKg5268+tV+zWI+POEoiQtIu9mzU+0m
u0aGltzw4+TNgbv0Z9cgH+LFhBcgWOMJQsNuXM36Y+wrkwJ/cRgtPZguJhkj13F6vWc1bTBeYFUK
gIWMXtFHqA+wb6L7h94NC4TxeFJjcKIeH8wP1krfv8ozpzUcdWaD35VWehIQqpRWfsXfDiyeb+yU
8SQgAvTaceYh/NhTuePWQ42CUaAgsOwWmuBkOtJJmheVKlkYsg3XV5pET++Y99F1GnIY750jvEow
VS0lqvpvohO4k8qr3VhEdXBET0O5LOadeDm6ei/+/k6HTjOPe6IG8Ykop+shSkeMYjjCKoCIxgXR
l5IeAAybkU0I4pkc/31y6uWKO/TeW3rlWc8nBZzdzyRYXvf9UGcm4lhyPmCokMt6YyzEfWvNg1ZP
+jNtfgwOdZ6+wjd4i832TrdnTET4QKspUeDdZh60xkqMxYxm69Ex+ifi0EbvTp+d/rPLxKuqqMpK
DiY9c6k0lNpNyr/wChjNGSaEIloLPdtvxiTRcOq34LNQEJxLIeixRvvgfDgcSmBZhuNwVnL0g5cQ
cQEYDnHv2gEUXotRIAd+W6TJWcb/NA16swnIOCnwJMXKmvlOG3gnL8nloZbxaVKXzEKYE+7g9tg6
rb1qVPwcC81aHnmGRoBb6cdyk+uHp3cl3NZTfRvu1tOQlgmp3kgQj8lFOcR+buoHV9UITr1X/z+d
QnF0Nmtv/FkN+C2wdDWdNb8bqScszhhFoS2/j44OIQBU3Jye7S9+UG/TvmAU3vWgjJ3IqmkeO8fO
QnAUONlw3D7YF8AA9cuIXbHZIFcNGO1++5peIq35Vkf/v96JS8OcnQQHI7RAmZq0OCIdpQ+FlLBT
6jOQmK6aoBBgE67N6U0uKc9u2/ZHBtXlyOjjDHiHhEwbJZUi3EhG+GnDh+6Mc0m99+JNO4iC4Ev8
1AdrIbJSibosEBhJ7gXDeYLTlwmZmGYMmB1oD/f1Mk4zrWqGg6rmQgUmfe8oVlkYIqNBjkQfaCS7
RHx/ctaZcmzTokT6SznBlwDxdmXYlJmXHUeo7EAw4PHvU/hPj5w90d9B7Q9HSRAH4kLKCm2kS6EN
tHsZ5X1cPCISPPc9V1Z6aitg7kp7HF787AsuBdwSUzEd7k2+ru4dPFRhuj051iGLceWgutXOFKsN
31q+QW1jKPVxFXkAAJQIabRrIE0Vg/Y4oXHrCha6IWHJPZWpA1l4LVVzXfmFZBikvCHmx9/V8pj1
DDuP9CGbVRyuFovLc6bxYSfCpCSH3LXvhRPC7VjAGlKv/hecy4Nwo0SQIgZ4dJSS1epaCJ433+IM
2bQmJ+hCMrBxlgHAYaxFUmDlKJmpheGl6uoTTQabxg0l5Er2f210rYFs8RNbdfbp0uB9R+LQ2CZE
E7xTaQsRqbIDpj16gSy59FsJLK7qd0/iFIr+BvHuw11RgT+2uXPdHYbIvwc68iJ6m6UgND6v2wzn
cq/2i/c30GFc5/5/XeGIKnZeH8VZBhgKkLFdspSftqSFp1+OGIZrzDgQsKZ4Sz4VetTkuDiuzQY8
xDnDyete4eGnx09201ZaQ7YpzmVmqEQ6pUWB0kgyN9IwAGPjaA9DnokBYBeP8fcsZPXabsUG4ClK
wmGqKRmKAQsORu5KlBeBCx77TfIK0d6Y4jnnapRtKjSBg7z3U3Y+nYJcFV8BlbLBL9/xRsefdbrY
jVzAvbJ8+T5URLl5CDi+WmKUZgykGfbL0+3sCQ6b6iyMzt6ZYspFtBWS4qkgU6S22z1jPHo/C2gE
7WAlXWPT70CiZLoCslmjO5sVK5yWEHL4MFzIHUT17pfqA0YPWjV/qRVLH4F95Y1McFta7FRdnaO9
Lxqrsuw1FsW9zqQtmxboNymJvHLD/poiiBe3evyQp1L65EqwtzU2Dh0jWWzXEAH/8Ec9C7heO+eD
wBi1TxjTddQ+U8MDRDPPGQ1tRLFWPS1LGxIAYqz3jiOs1u5AwxpQU0fQi9jQDNZLfSUh/OPc+U6N
QbC30oK4m00CMKeYmS4LFYGTnaKxy1QYnZohHzsYlNmGhmlh6Err9Og0JvkgicoAiKSgJNQdWLo0
3iFsvOGFjtBtXBsu3CyfU/7IT8wPg1prLzs2n2dh+iP1Cb4p5M6meHpGJsfUfH9WgoQDDs6s3ctx
q80GXTJHaR0fz8HTE6x4J320keSps0/8sYiCxcZPqjbDwWCOPE/V1JOE0NY9iPpTxTz01Qv5hbxc
Gskq26qfkTZRQZeOL0KWAyoMzfAfQ7bw9O1FDbK4H6oRUkg8alBNcssxTTcEfLd7TGKzoYvvKoTp
BkdwDQdkDszBg+N3dm8YyjK6oa8tiSCv/kug72cxBE7ilLpd92I4UqD5zn7+Il2PMbSop1MWciva
AdbucTBKf42nrO/B+ELJ/8W3zlYr4ZxV+qCNWewl/7kBmwqR+d2bvxUk43yYyaWRsP4/difBg9U6
qe+9YIdzvn1M6DB/G8s37Z+43HiU/aKZEOzdX4H9qsL77j0ieINRepi/bwQYLTaWAfFtUg4nXs8/
gRrXaNUEHAfHphlkagJPpxUdHP1aMGLgRxXaWg0HfNsE3bXJNCaB0nnBStBtADqLDb5OCUonjx+o
u7IpX9dvSzVwrgiJCrF7Dq3LRCdx9QTiGscZTypw1hYUAe2Abmq3+o/Nd/W0dNvhvjjiUDz4Uth5
c3OlLa91kE8TQhmYQPugdFO5U4FeXrdh/e9RiwQYJpHHg05JFNYIBTn44820LpJ9M6HH0U6rYryb
wCoQtOio0KYpKNU3v4riHIB+7j4aRy3ui95WHlo60Z6f44aY2ZhWCAJTmUIvBVKzbQMLS0uZO+AZ
GGzZPomr6qUu3h9wt3uCpOvHkrN0BwKNZsu9guPNgdeOywPey8BCyeZm9i43iECANVKsRH5SJyH3
KV6fL3rV6rXvddnZ1mITzq0CysWPBEuN7HzKakn4I1NdTuV9Oquv2IUZuKjV9G8Qnwa+WRUDHGV+
wsbP/J2l8su8qHWZZeJhmLZO9QaARzLDE6fPXiZ6pg0n6qJ3LNz4QbqaVndBBFmJlPz+j67Fme/J
M+Apl4o/d4FNw2eU77g1a0WC2poyr0J9wCdQmzxNCiYj0F7EP1WYhIPnp6izL3DaAaPty4hS9Rnr
NOtyIby32Nq9YXPDlrK5OGMOfNa0A+DlC9uTC4nCqnQe67+Unc1f9kT8AfOkKrXbGEJ1uM4uq7eQ
WGJdZunna2sobu7Q2tgx4mxfiqaqG67Grw4uIU1GqGNSQBntsMKs23EwzGeUD+rGMvUtkGmwEJeP
cW0A4wd1n+Q80bLFuJOLCQH7OCuyeb65+os+jNZTNK5TpVWZDXc8qv8TxgasbddMZHunGMx/h1Z7
r9HiGPkCACzRorARaFpNM4+IIypXe3q4ZHxBEPE0gV33jX0txiiohFUYIgscjEj3HiPEeHqVrK+q
x7L/UFwSyrAhTLswLkFbWe8Jw3xE607N47wzPzqnNweUU0GbSc/4aJ5SgDa/dmNqVppZrrEyK/tg
vksApy4QcG9hqY684/HWYn8d/tOQibga/hhTv3RIb9+z1lUZYKNm+2KXRMfzJRJAFxv3m7YwZeID
qcbUKlQXA9GGleJNAPe+7s+BPBIdczOPgf/VqsJkZ9QvfMy+tAQ5JiG/foTExuDNUOWH97GGxHQT
yYAojVflmCZTBedq6m6tQL8a2NANXPhs/9O63vHn8nh4kXNgs4YAOZ6C3WyWJef4JR/UWReUyuVb
JBgEdV9JQXrrWFEZ5rrqSLKQ6QbKRBYkv6+Kzx7Z3cdRb+A1J15+leg8JbfM+scIC+d7f1UfD3sh
Ze3qRYzIsa8Hk4zy8mkMc8IOvPGGLlkZKhNt5Y6VAFG6KDYsDfKUOtsVBYgXLGbIg1xzW+gBU77t
MYnxSAN5uwqQLu4bwSTVIZKVrM5FjLt/v5nQ77JdNJrNc3/8ym5P5L33BXq5kr0poiMpRiaVZQ8k
S8rmonOrXnG+G5+imMZ+V8hy8YsDD3fyOgYHcHnyZ6Kuz46PDeTe0fu+gGUv8JjjJFfhZTDWVraZ
Y1q9gkiCS7aN6gEHAyoKmTtN0w70bUs/LI90rQWbr0f19kmr1+681uqP+oj7flScqbQjlw9oO5vu
9Ku+rs3c11lRaqhnw8GisladayE9hBnTxdWs4ui4DgE0cwL0cef0wTwJOMkgx9tKsZAXch4gAzNB
JPPp8XGsxkoB1nItHVyBMRK4z3nH7xp0VLin51I/H8oFZKW5z/tygdOByP+Bno3AUFFkhMVq+9mT
v3OpgihmSUZsMkEfznkdOZ6TEOFNmKCDjrjCknHBf00JWEwZYaCYfz2ogekxnwtaTL2fK7V3acGS
//hOSnRdCVLWVZRZpxvgJFRGSpshfqxjRXN1DK5MAhHXFmjv9sk1OMrdKG34fnp5Nd7hHJ7x3rV6
+7HOxT0QABMNGq062fkOxJu3SOFBbEJRMXd0dIt90xrS7ARbIeN/GAs+sTgAlXQWyoTAY+n8oxui
XnKabcNzL7RDpUy0dCwc3pBcq3u5JfJIe40Zy2pmT+iWNWL0ppxw8gT7jYTFNNQ8wtyqAAbE3gP/
OMovTTkHmGFGFz77aqObgnDbX/sfqKIV/ZUlo5TaZl7WQLvyOz3fwivnXo0z1wmrL7wTQYoVIV8/
N+7M4K4iRf3Xiwo6MkYltIm4OS1+GCdItVVv/+1Xi3qzKu/psB4nrAxuwhWJaGUVh/WvTKL7vsRB
h07gpc+AwjwloSYMoQ/SBMZ9VLMMEF4nTppZaetGui/SnZwvq/qUXvKdw5ZE8XgRW4iiLTpeE4k3
f7AvjuTqE78Ao+NEwBY0ya/yU+6C59FwmqX0RvHYBtBnlDnn8OJU6HSmz9ql4gHvpkuuXm3S/IHK
s8/cGWc9c+n+tGf+JQFZwjrKV2TTobESnrE0hYPk4QIYX75VkxgIsxKr25KzuDj6tSZC6XLoWU7N
+5SzbMuHxlWVrbbZdBlRa5oari3MzxC4+W0fsMlZINn2y0ZBJ3qvFkKFkvbxr2Wl51D9hKqHvj0S
MLe5VQG7b1dpTySH+LrgHRetnIhpyI5E+J00IIrYrZ5qb2vb/D9k3M9kk1AZ9ecEt+qKDY/thGey
NrflQJ1cibOgU8s6B/7vuCZEjfwtxTelsBY44xDJXQ0bkassvz6S1nXX5OohLcq+OQmsm8hHcEcc
DtwDhJF8OF9nKQbifoQ1g9wop+7hW3P6atBDheaPq5KtrVsgis6SodMAQCzPK8QPbMPfedEwCKFv
okU03dd5ysSPUwE4Q/4GZP0Y6IPZHj+4axcNPe5Q/n4dwqKfZw+PL+64lpVE399W2hyQiCS5YMlI
KHByRuHqaUJrpNQRZg/PehuuZ0vlVu156yGnU7w6hXhkWy8Qe/7dlGQfx0OITjfheborssLoCRQK
XY5XnhYTOgg86cluQQjGTpHQBWq4qVQVtfmVX/AgswJ19Qsfs/x89vF5H7Ia2/3cfuNrNDPmRlfd
v126GXgrcm0cjw6nhrDeavx4DDzFh62kCJEu4MV5esrU8r1AiFKtMPtKd/eD+IGhK/Y+a31hG+xG
TCRKhVqE+5xLPXkPu1YH0Cf9mtgM2yYIpeIU00dx0HKnxYi7dkr9eUQpg35Jue5CfmZJ1n5xHRTv
cl5CmyNe8IMMzl13penvwXLPiFCyo7mtdz3mWIPsaynYEd9zDvmOBcelcuiWC0M2WFwO+zEs7vup
E7Ntq9Z3MwbvNQybRzEfkXxk2zIa0NLVhpkJAVls3ubzpYw1CWTR8TZ4WDfaS0TI7TFrT8GvrCIJ
9o0Wi+dvY9Bh8K0Dd71kgdi86BiB+vcWiQXgm0RstTL+FSiwXwaGClvA3TR170njHfVZlPq2DfJd
XibjGCRRBekW3lrRAiIyVRyGTNMwL64OMz3rIEc2RiLhTTh55IRUTM1YL03ubqAlQKI38iZxL8YW
LiD5ThPofYUKluqDKkcAAVVx4Ku2Y/bGtQHUNgB4RbHubF6UrwygzyzeUA5hdJHAj4xGu+bK5N7/
ESwaweBFBxI5y755tRwGNRG7OuXq/wAdZM/9fedD4yG+q8Liq04/VxKnkzfLwbzVNbQNagS8Uom+
CxP3edkL7uLqSv1+EfFJl8dsEOaZ8vek/zN6lxSb5n8/1lj2N6YtGhrgwj+z5oDj+tHAJ1WdLzK9
9ScvCehYvPSg3p6oC0aw3u+2imxgPSJ+KPH02KnBAq91rgU+N9z11Gs6cTqWw6wIusaw6HV6nCvZ
2QUofBmFK/Ei/+sMP5NOTb9GHX509C1ktpf5VQ40ZmI83pOwTdj1MzsZo5weOcGnokcXjC6L21aB
zDIXffDkiictA1YSv4mI3GRRLF23fapLOpfa1YN5WzwbyCnfNqBHjoAJrtXf8iSEob0DTlBxee03
27WL1nw+ywVBYAy4+zMkMLAT1TLOLKfo50y6hQzPmcmhB6pXQ5D0eZKaM097CzAcmMJPhxQbuG6g
wqWe1ZQ/Zl4guh6JHW/PgpSJH64gXQlMGQ3vXd/878jYm+D6f+Cuq8WQbsM2+f2V/+wbvA7sIQtg
vCzpT0BC4AwxupIypUO/PiHAFgUSO8qT8D+mlGGY+c4n0Zhp8LTjFtpo0CF5/OWyiA2eghkBTrlZ
q7zQclad/C3iqJZ133cNfgtFxDm02/RYviIbF/coBlYkZgn4YKJs1eJdcpYxg22wd46eodsQjbfp
wFcCPp+OXos1U+z6NqF00vjKodWjHURlKLDi1rAfQxYQGTjcRpA7fngs4Fqci5OAWcjzf4DHRmLe
ZZh2rOAbRixwawJ2uajr6e2NT8Skte8djHNVsMONOyRX8ZHO9oT0+KZm0umXiftpH82RmEWfOBOo
FSLm1TUjPGkCuqZrm71yS2mbmSiL4GODX/ckwjUUSrdl73ICm0Ou6/TfJo16T9MdJGHvdVGtanoo
7EgRP50os5jYSs1YrML9neyeVZvPHLlIchTngI1xgNtzoJfFzn9qktWimvvZ1FRGnrviLoHoH/LX
1Z+BYqzxvhl/9hZO9iyK+hqXaE5VmUNj+G0sd/OQYmVXN50GGtiPYvYggBOwFtAqkUfDaZK61ATz
istPjppbObYH4nKU/MoHibT01Qm4uuC/vZ+wYBXVG5KW0WeXXoDrVZhpZ53X+gMNGFKyjnxO0D87
ClfvHnfhmsomuQDoX/a+4f4/lbInDvSR5FQbYl4AI21CdSwh6943iMR137mmrzFyiF693SrWPIXT
NQV5/J1bJyMtcUbZlzvQp120V0RkP5yGtleLKFmSMOs/uFVggMO1/WtXv5O4s4YmxJqKPbFu/Ns8
7FDUAz1aycZqUEh8ZET7NxJJj0El82NEU5HyvoS6X+FMNWgHLDL5cbP2qmzYId/zQ77W/a799ftN
tieM3HMWKRUOPzsxEYWZB9Vww3v+7F7P14lY06n/3hQ2fMAzANqFbDg92XEIeXwSqUnW4XXjoDFv
SaGsCEdVrsUiuIBPA81UH+AyoMEN5qFN0ON8rfefDK/RwR2N0+iYs7py50HLGN5sqZXkFJjaHLpG
ZzBYvw/Z2VlSdSblVGzsdfpQ/BEE2eIh1BmVEU6ymfL7bUSHWAC9jCs270eO+Um4raVR794XseT4
ee8Bb4hZgbxy73a4rs2j2oVN8MCbctvUHZ+RsfGxGW1M7NL2a2Vf6y8Q5PibZOcznGPsfanurlhL
2J7hbfmctF5bLjbG6EDt+skp+Vq6bGHlKYsiCdKzmzYRUZ6S2e+1/tC1bOuSWmPOltowOfMvTWv2
yV1ysXLO6COUjB8IkD/otJGABlByHs2a/Obp9Sk43KuSQRbR3+BKK6Muk9Vq5OX3iAvQwilt3hPx
WAxpm+UIFPVzARw7Uq/q+y3/hVV51jGAQCVkQF2myY0oiNibGWtJSQCF9e5DCtCQ6yZOLEYVLRxR
8kUZPRmJsW07B6QNosfLSgYpx6nMu2SRjY2inB9JagSH6EIlSClcr1aIl4hPJMnQivz65XesXERo
ubRxROWJyCsy5eSMOvAQM2Rc6NC9/05n3DDgTkeVObL6fWkj+P17vsBd3VEO3MUTsr9bmMoQWpDm
b40aGkLpFUHJ7K/9325u8LprGRFhf6nmQwBfy9jtu8mr4iehGJOkTNgHDCDQB44EKnMNgdygcBWb
ONaVTx9fVvLl9CxSVE+9C4tbnIikBDw9HvYq2I17jNUKcBhVePsOyja1lemWRQtrNC6nwgv8poPs
8pl+5rHTo8O6+MKi7f4ga9SVgmMoQAInMdaE3qqKF0/zzEhfjnolk7norboKZdOloClLtgpTbvgP
cxJsyBKHUxHGn0WsbnQc/Er5nj0erMPh1CLzMKPFJiR+oi97Lt/d2SJw7xyra4bzhQtqfHtLbNZ1
3bvjo+OXlNng+7Ud5b94+AICIJFtUGYg62yqT+LgRBLE8pXdyLJ8VTsjGjbx8prLlEcn/A2s0hdi
WaCO7YbIJiCTX3yI+yjVZIiXNX6ev5lNDu48QoPzbVOKfeehASLQKmc5diDWtcCgd1EQ3z6jtfar
JV2T+y2v7zI66egRVvyTdVefZW2DUZta+KX5/m/NV9DCF/8zwgajgY5Ysl84he+fHgRMRUUNMm1N
oR2VJpjpKoYgLqhXCZEaJPLDHSoU5nNLgWd24htmvQevCQeETqi6SHfbvyucrXkgO9Wz3u1GRY0m
iQDGvgF86Zmp5AwcDYgsM3GMrS+dc6c9l5SJq1hkUoSniypxcz4pjByvtYFjr9tsmLZsv4MUhGY5
kqASQDJMRNN2+JEKWEjl8Bq6a+J5ebEn0TXHbTXB8lZU7RAyX88OyxysCg139vy85k3iTT2aONfF
xpQBPCxF9fkSC+F8KRAV3V6r07i7AFSwHInhKIyimWcpdL8XbGiYlDQFeZnTDkTJ1LN/AH6ybONy
kI9Os2TsuKwVehlaRh7Z7LF4aGh/aVeTlEvd+me7i3wHOws+217bwCWFi4dBfUkR8TGqvZfjqovR
wPrPsN8jC9aCMQkWuCzbyUmXjRF/GJUkOmQtNOjmuZ2r0Iq8G8ByNiAd4kvN6LGvRLzGp6BSmFHB
wNvQcGQ7+rDLxUOz8YEdAlA2V+JcV/NsMh1TYnvSLt9IZJCAfTBqozMTpaHLFRbPYWkQwmpWtqS/
nGYo/nPNX5yexCVdDWBO+zdXet6z5VXie2ck2QrhyN7HbFixD4wJuPMoo7H1HKhTgQ7uBi2GyHNA
132NDj2ypdygdTCiVJjV7RsPBfWpLAEvhGku2hmqXWeW+dzRo/tWlC6ODkvKR2lGApIw6IoOOgKo
GQ8lLdU+ztxiSNdBwJIy1cUZaNSCoWPo8vxzs0xnZPeCXVvSlMvmElm81+7JMj9B13k8aKnnz4u7
bedpV89SHML4a8wwCRc+lRGnOwagYR4ZcdCMfalYKxUqOriPXI0KLVtPj+JDNcOd6FIY18W5JGKm
wGotSfojb02ptUcSV9PjI+MTeH3No6T3hZHC1c5Ni5pH1VmpeQCIGeKu2A5CcUugIRmjhoBiulqM
8QEZ4k3Ti7rDGYxvbuCT2crrgjRtpildrL6bULq4FXZibB7b/jo8hxygBHo2Y432/4SanGgjFYJu
srq5MBwhlaUWjdpNjfSm1hs4ckk1osMnzUgIMtnRL5nnBu1yU+DN7Jny48+xLB2xjVGjwF0gO6u8
o0S03TikvTq+NoEB7q2Nz13HaX+ycpsRBFroSdaY0DAVXYvGLfoQGCaHB1jXeDvjTUvZX8Nppwc7
SgzhXcOmsOfnQrknMqBEmMt6JMixiV3VQA3qfIFEODDNAYY106IzXkTu85YFNVeJDUQ66d2sAjfl
JtKCUUJuY0pLPILOoRZr93P24/aZFcLdKtURd6hkWIuA5YtMlvaDXj3xzAGn0OonhBTFmyvM1Qh4
+qePthFN4URv0w3mMaoydgNh4ShIv/T3PVqV0xOcz6uC2/y9YT1sra8SHug8JRfkhRaTPokRUx/y
1nsE8eWicSLPO04xxIO1KeaJeDEXZMrE3GtC4HI17qZkcrrE7QY0jrAibkNR31dwWrUnZESMTDn3
aV3CJ8nT48WMDLwxIvsnO0HNE8vNZCNW61GrfM8wD0q5vOVIOldr6epOp0YZYItSmo2zLK7ixhs/
Tvxzjlr88pkq0P28jhx7uEGCuvXJ7HAL8DcUd9IneOy3QF68KypHViX0w9LXd3gOXCdvB2HCf7t9
G5Hou0Z6rRgUzWrlpzLqow2WSWyEMUaP6+dUTF/jAzC7ZMxub87qaPcZdi1pI+yN2O+fyafHuTY3
x4T6o3+rNG+YQpd7eSdVhLDmoXdlDclPmOieqmAZULkyAIgyyFuaziTWmUVeHsUeteeGF2CbZk6/
ORs+ZERJs5xN5LXk/L+ure5VLIN5uA1Wngo9OQx0CHR9sH9917haq+gdoCFanYo8vLneW76CC0TY
rYkz885edwZhe+4gq+RTzDJznapOySeewV8w/TYR2qM7Gncn8XCadINHGNCY+ByUJRapXiQTP6qy
EfS2UzqSWLKP1tRLT/5QtZm8cHxV4G0uym5QX2Ziw0+gIVR7mzBAi64V4iMQyKgXHVbKNwQKStJw
UGR1Y+f6W3w+j71yTMLDtocyPenIe8JuUKVYu22S+oKGMUOw9MA7qiDqutInI+ZocD9orhPXBkFC
LWYqctGdWq+mmr5XOEZSMkSGCDIGDafNlybSQUzZNo+2cvTkQDh5hbXlHffasbDt+AM/h19S8K55
oLvLAZuT8jevoAs5vrBpfLojSbgdzeZPvnUOfpI5xgKVhKbgH/5zvyWTpV3L1537H7iBJVRRqVHr
9W69hZvxXkiqNZ3P/+o6jDc3rZQNCqiwt2Ng8oqx5LaAIityIQ4TzpjhaciwbmB+maRYVC7OA9uh
xCeeaYOjhmEYqT8lz9JScS8jVT9ElEvJVsAvYOcB+ZZKNZnuUoaIFMmfHOWeoel703Ds40E7cSAd
hN1Rt9oMdk1CgWnze0zBjWWVQr0t21oZjKqab5O3/HmTMPvuqwnYbDZBIpfIYWkxX0v+8x8Wwsv4
jZzutRSfei+1q9J2IHRFYDKN05n7DGDDFTumDuf4Wtd91Fp2YYbBnRILuNW7XQE2DCnL+Zba1GqJ
ECZVpr3AXw0IIqdjm2ZehB+UdvWQoGoqvh6JTh3WcPEklSdu/QzwGZgoTRHE3RCE7+7uI11NR6CN
VYztQxEu3QD4VIXQS2cbvdjNQSTlZxMabAotJNwPvvAXcrWX568V9QndVXm5nXAi02S5NeTqtU0y
K+bcdMUDmGlagFMSjhEIOTwwCkfkfA6H0hPrsEbHLuGFgt5uuZe9Fvd+fJ7jtWAoM4H+Bgvpep03
mGSWWD5f5MKWWbN75R8UuEG1f9WgwdVw3/byp0MCJGybhb4nUZgCtqG9X/VxeUVsPlpvSctMgfan
KKklQXvlJkafML4B6gd5F4V9UiKUic1rMS6ZeYphcHgV4FezY9R0iYQbiIWqDD/ARmbtiW5uIguI
3JgStYELL76NP8bekeK+zd9/zUq+7yuSzHw+ZSbITiywb4wcOQav5Dq/eXIKrFOw44SEyiAxlDjh
A9kpWEyk7OQTGEl6bg9xmf3Ly/jjZwHgT1VGhPuTKe6N/JdEQVzrewG/CG2tkVgsw+nTU4RUxBTp
GGRrqsxI6nTVFW+u3eUcyGrnNC2LdSoHjduTAQI00Ij9awLJ3sRywSZU/pmFMXWdicM9ArcqOMBu
VMkiWTgG/+PHCEQj9Vez6AMbeE7dri8xokLrFksaXHRR9yyGTf7DHjMoNxF1QdtwDSU1ydX3dxCX
Ur8RpB+zVj9sEtYG101DTnJcAQlTYTbbU/Y/g57JvDFT4ckY7iOY11PwzLftmkyHG3oljW1nWYgj
vPutFzzEI0DrSLfCUtOfLaBkc6CImXFvQehlHLGZE8PQG8DKvNoacdvMkODgDEingIL4ErQM2ZPz
Fp5/6dbt58wOjQ8i2vtWB+sBYq6XLGT/8p3VEN98jNV1WSEXjutqjesG9YjHkn1ZXa1bJyq6rxIJ
GF7cjWsucSgUfTAfjEsaIxfxtckojb8+yeClQwRNYadEfl++UErhtywaOoYXkAcpQ+5GCW6BHAwN
ACmu/3Qp6oIqq2cZwAKm7vKx8F/0ZAZnfjpwbNwLobB0IJO7d8UEDqVwndeV1ENW9lbVYUkg4ud/
OVw9xTpvg0cx3w+k0THBXqAYytNiIc4Hs+Nu8i0vn+dFdLgdHz76RTSPgwvnSFOcvYazZNXAUKIx
RCtTUHwyLD2a+YlN5S3705JZfmO1ZEDD2N/NTH22O+7SpoI0yizCE1Kg5VvVFWsqo+5jsbcbpkOw
Tq6WJwM7+eVo3KVKqnHtMJIssk2KFRqtry3RFvxMaofCX/G/by8Qj1IRg/SDjI7CDoWtgbhNReer
+y5oQR3WVm7XEyXm9zQqyyC/MlO0E1/b+8b4F9XXOe+7WB7xJreB54FoJvat0SmGfQzWVUCTNuQs
THqgTra58M2d9/MULCG9KdLCf85FQ65lIcdgCFC0MSRJvVrm9L4FWdeImU0yBSQ1nv7662nHlRdx
QP2s163aPeHTrtS3zvm4atpGjbkdVaY3oMML9Eq2Q+915N0UnyxwpMm3aC3ahX6qL0pDjN66kE4j
AkgFEjc7bqF9tGqwKHtI1PQ6oVBlitY40bt2NSFNlFAoPIgLDPYFwBf88DkJ/q/MxJHg9ZLNz/GH
xj1izzRCzM1B825mVSndgW9DJNUpcLDuu1zQWb2wmH3KK/TVis2JzkQmgXpi5JYfepREmIGwhFTW
pIDG3PT9xYa6kUPs+YraXNE2ZprSSgdYquEoVaYNitafPVAqrquJ/z4wZiSvhwqjjV0bDgT5ItuV
Ry+EUgKZJ/VI0b9r88iI+7hV7k59RQdf6up9HIaCt4NNOiMFuMMkM9l6IS+cBNGK8l8vbpWWg0nI
mG+fZpFQey8XBudV0z8dUmaz0sqD90MQYBq6lUUltkkMfoytk7OjltpHVet9L9ZPqBKsN1lTJ8Qg
IThBRA18aCZBeES7rEgNMwZCzxG7wWgZ61Nz+ekHOqRnHB2trGqd4hyXopw5FTYsUG4biJ/4jEM/
6zNpihREcvlewGzPP7vASSK5z9bQ+2dxpqYD8A89Efc2us3tYvd0ol5qni8USadlCKJl8CysaR1t
77IuU7v+zD0XXdUh53WQHh+63nJrFaWzZJhotXXfZlw7Oj+cUaJ9k1yKdMz9m8rlyRZj/cuuc2sD
fiZKhES9I55KmfX1cU+SaiPHWCaeS6p1VYwtz3Ird9a3uwppVrpUey5aYGno+JV5d3puo0m3gAvv
TGVNIUq2/wa17nUESu3bHnc4XYprAs7wzEv4dJELJsH6Wjukn3zvqDVrL058TbnvPQHktThJZ2rw
9W78LvvYIZD9pr6RfQv62kWXBryldqV11faxx8xX0bo6dh2IdZ6sHg9e5qK7azMQVi4r+rBnWDkK
2tC9Js7Pg0ez+Cp24P1rrygDCnGf+fmcOx0R2vL1Vd3K7qwBAwWuL/1j6mIXMkWR/L3z76SLZI08
8FtzQIA89IhQTR+GZcLIQQf628FpJVkNuLDCPBJAW3Wj1Ak4hZzIAMbCp3Qe/xEP4EuEJ+6pM9q+
ARYmgyh4rYE6IwNHkfGQCDy10NQ8T11Cdieul/wKNJV2fl4aQbJQU4dtfkOfcNm2Gyui9Pr8dBni
SrB4Ch8f6OfZdNvNtbjBt3d7QnqYZ1aWcCg5y6b4kIb/bw2I+fKtRc5OkVFjBEROCCO1o1/wOD3d
jSLTQoaFY3QNs8bHTFe1qMllXM4u5xf2HdbJyeRQ/SuwxxuNgZItu7bjVTegl0RIp9A4QcInPzM1
LzkQksX62C6GYKo/FziZAMeQj/fgjjAv6NjQdQ34RBzJ9r1OkzV/uYXtLdHK/Ttzvw6RF9oFsELg
OQjUy5BQQAFxlsWbQIMLteFuxMy7AD8xMjHQZ9BjDfEJAoTvUfb0OIHZV4IL+qSkTeD3TkyPGPsZ
5T0qt+Mtc2XaIou3c8nW4+K59MPpEZmYbnw8TssGiaohjAldWfJ3gV9L66YtZJEZMkPSO/xRjlKC
6ZayDOrhD4ZeLqymbjnkqgWo8z7cAyyp+/lDfk5bfrFChVt19xbqbqUi0aNGQe4CdFnpsKeZ/RMw
nLiZzrvxN0Mn79Q+qiq9xwW0W+XcO7/Gn59RWTG8jNDvo4VTsS5mdhN+sWjpe1JoXyKuqKu8AK4m
P27Sv8QmJn60jVT51dN13y7bMe3rsHLg0uxC/PKDp2o2qN7PC3xvtaOhkCyk6oBp4wQvSb47CBsw
dXTTzzYNlUDIEBey04VPKEYV8XggRWVk5QkPELx38HDPb7AMoO0TgwBFhIa4WzsgglkuBVo8yMIq
w+WpinT6l3Ig7629/vI0ig6wipf585zexwBypsAi/dmVt8R2cvqY0X8Di70fmymy46iuc/FKHBmS
w0mv0ZKUGoMim8h5qzt0G+sZ+iFlXnejMo9YdCADVUSE5zk8+G9Gsk77QlqMuWOPdcVfQJVTBzBR
mxLoPfk0ij6d6QU9BAcoJC0ogHvSOOCHnQpycivPh/CkFRpzKlKxdi9A2qleWVYignL0zn7rmVFC
27/xquM5xEYAj5n9NFjD5u+t9WwMv7o8alRhm5UwCU4AgGxQwNW2GuHuqhmfAgJwUUv9pWB8oIZv
JHY695ASdqPPlnzSZ8g1v+pxxpwqUdqqXL83YhXXNXTStrqyXSwgHhtQn+NskqjcGe9TkQsPKwuE
Y3ido56WsN7cKsM6NNxtko7N4eD1ZbfpaP3TrjnDvUlpdqQ4kteNXvMSzA7Lo+Uovsk+s3WME9/P
1DrSXIdx+0Yw0OPZHCOQhrUaCDgCLZ9Tq0ef3mmzfru8EMXuWnxF+aiWWUtyLQPU2pCLNmnYWAej
0TAAZbW6hIhqfCbFUnODaex8bgenJ2GYk8bEhAPU8ZLW3QhzJspD+0VVmI6EirnXIer0pXjNVF+K
ro0u9Mau7yBnmLUB188acRVr8CeK+ZmUHmMPJ9zATLRUy5xbzjvNWLZ+uMURgIhIKnDy98rR28ZS
/gLaZRr3sVFK84BS0CpY3XdmUv2ZQMy6ETPPz93Kufug5mX1y+vyM4eSpX4EOg4K/DjjS9B9Jygh
jEst65cy7GI7nX4A1tHn/JVTCM899Z1ENhyz7HHHBreG/ZrhFL7qOgYdycGohLnIju0cUMDwtLZq
ipbGzds2WsG4wqwrK6HiVh805167h5HOXPQTgpAL/riRIdqxW8xJLkq0T+E6w3ZgF48pb6i6FCS+
oyJekg5jWnhExZrHZSBynp1JTZuvH+mELOTO0irZRm4lIcrYIcKD4LqoaVOK0BY/1W7/Mp3swfq+
Sgj4eLD2GBACdctvhCs5bnsu0znc11kMW0zOxQg5SphYCxIQ9nfhH4iO2BHCH2piuOQN/U6RwJyH
X0D+g08KIEAUBY/3T4Mdy+KjnXKaqrz/ijihM0ZI7W4rG25AGxCNjmrn+3JmUbJ8DjF7JIAiPOwN
2AYqFvnZMt7kivK6M8Gt7nKPaWAd4cFmmx3IJ1RkdyxEXCd7bs+5aRuGGVG8DdY5AXGfxa/tyld4
tKt5tqC2YUrhYEvKvkQxrLUaqBeBcsCGKks+utojnQPaumZf7Hh4gO6CbckUbteAH1mzWx0llxbN
GI5IWrF/M4O8S4CemOtDIvZgEz3NjBQ+IUAl9Z3LoiHi9gpi7TR/dirTRRtVI8QJn24F8p9Sw1qO
ThWKQLPKg5wQFGjdcwkA9fD62Z1cHn+euYQ0BsbYZarw0bezi3lfvwEF29ctwvGBrC5cpv4vRw9t
liWdzfXQkDhnIaU4+PKpY2hGUwyRBHzf/uUcK1OCWBrBSbOjbV5+PuNLMD75xsifVvdk/P9hyqyq
qPgfUBq4y3Jl46im2kXTfpuY+CXAxTt9DZPoLysrgx7VsqAKQvDHYRO4URtbpL/ITTKCflEGhwnZ
cp3bKDrh8MsJIF6f9Ha/rtQAyRI+og+ZolwOu/STk0ifT87QsHwzHYDZCUoLYtahDGSUFjzAaK4h
qup1VIrH92x5ZGzhdiaRuo0mx7JgOsA/XUFh/F+mTxahgoOkcFnE4/OJi8VzrwEovbpHz/DUfNzr
HTqdlt1p+hSg/cybteek79KY+83OepY41t9lzLYwcQI1DkL+m8u67wjUah5nPNJCK0NKvORtRrDc
18nILi7OIawnZSKyCuTIt3eOcDA+Qd8EiXhpHJlcvjE/5ElTH9KncJsUiycrYuXpR9yKYiGugvMB
l3E/z3maDoiuLCcYUx1sBKKeHOJsX+bTP7Q0Z2JsMGo+4N+zvX+hvFRH1SqJK/EDlVnKIN4Eiphw
/ke5EAci7cHHNI9APqZoCl/dnCzkCmffHfL/29zuWebMDGjjFxWmSm2T7Ww0xxtFGmEgUl8Xm3VI
PeFQ/PZqrD98eGWeujWxP+o5dr0TynpgsXhPw9WoQbKFSPH8VPgSPQxQu79Xyxzu17p7ME/g6JCM
IJBcqkcUcnZUBkA8kMn7nAGmJStNIxuAlWP0fxSvA1oD/2KgV8TA02kGjM36+QBEa43oKLMf/bJA
vwc7YXFLhLM/jsvBZdVTlmsvsUX8S3j+FhEmXK/D50nc6wABhndrUOusL2WNaVSDlxNIyt7Vt4F5
xxVo+W5GAJjQlzsiOSq/VytWIYUZsmanbX01+QpxJBvYGRNvwolQuu606FnyCuhBTEiH6IrhNDat
K90Du8G9h3lGZvpXxL88YwOYW09xO8PZ9qgFRwFcKjbVJjqXgeTQfG0tE0gCWyOmR+FQWJWTzIeM
0f5o39Lmn/YKPMB40oBMgWc9EYl/wbynTmCSes7bLF/mp2cEovQMuk9LNoEYyMJZf7I3HledXQFi
5V9Krt33GVedROlDWh9324HBsWjwqVHA+Y2MRasr3RIdP0B3aLtCZgCb7/xb1MiLOWN5+w0bOdF3
53iBYi8vEAK82vfQrC1txMfEhcx9xT3Bv4JCM4ONVMr1vszwTbw/x/Q19NzKXx9V9Xv+TIK31mPS
6tN3LVvRBMX7+B5/b1uz2NoBxTnm0fxPtMq4AJMx94mx38gYn5cXcI0unMQ2EiNe/0LCZXZmRJFA
X74CDqXp/jUlkqNQurderG394h/AZ4O2sM9fgmV4IHSMq+4hlD1+AqmMR2+YR5z/WnjEfg4SWK5D
pWWAVLzApKcXarvJYjeFCU+m2Yg6wcZ2Mkqt4yyP5tasBp7hElSXkH2Zw3465wfRbqwT1e1l8I5h
qi3WYH/0yzIIrKiNxONkG5oInb3VXUwc4mjDP1GaQAUil2/hufQ8gykbqeqmk362/p4erjzObstW
INPjgtU0m80ZDssql7SJBeKJCxzRviDffe0ziu69wjv96hnja7/TcRh6d0ElJFssbyOYZRQ37HZ5
VDoQXYPeImXxnF5zJy3BGgTlYsjd8Xik61p5x9jbIBLMCzQgWvIAPkS4qv5DjE+P7bp3L94k4nld
A+CfHsNzyx1Knjsp+bnxdVYMYqPS3GweLt8WmP0d8Ld8Xy6Vy3GQTalUWHPheySnAMrvdm9MqCHK
yofOy4W1J5VIpCT0pNUXs7j88PO6Ns6JRpnRGLfiNBFY4UH1fgpSLrUZmOKOLBqOSMXVG6r+ByOH
ib4o6IDlQhBXAO07xAVgSpA7+YzUReD1sc5qu2Pxihh7p1lNV83B2Wy42LZSROzmBF97SIA9l2jq
7zcvPMgo0uCxeAB1x5AmU16kpqqDR/6gytMlpJh+drvGVL+TEyeakM6QI8Zfa3tt4w3tAqNvX5iu
z/iQuc57pxqnzQVAbxJ4wJTKf9tVkFsUeAn0cTMX3uj4ZVErbL4PdyYBeb/up9WDE1iS8Pe04l0I
1emIX++/G38xA0bmmZT61qGSyZPYwS74TpXNuFaBq63L9gB9jxf+15Iel9ssWuq6H4elsjZup4u4
Vs6qSdcw+SPstPM+wgr0EcTddQ8suOrZ4rYSv4sNKSH6PP6Hb432yHkOMdh8tJY+pUGstfFYJ5sK
C/N0plV5Tv2ARqPBeHEav8qI+Z+AwuBxaRr8w1i+g/za/gNpTVZBGxbpMVfSh5d2NiXnyvqp6HwN
khYWgnnbh26qRn11l0MqCwWBv85DuO9ezmxLy+UmCMLGWoIMIbNm1ZeW06MAX2An42TZcKWr2UqK
DEx3qlDeaklQq7jd9sz2DoP5SrVa/+wRBgn98ieAueCSnHZypO7giI6jpGgN5GmKi0X/Qzcy4Axb
+oKwm/+WFIzl/JJI9Nt70kuXwEfeaR+NPgjlf1mIihItPEd75pklkt8ru0GdtPMOkJCHrYBHqQOw
JkpjsDUJ22ArHqoZ43DbK+4KF/2QxxbFxegCXsgx9foGoSfBOjN66fZBcSX9AYd5i6+5ZzMzgodZ
rr4XfpfY+lHp5drTBk+Z02lPCwRiBKWZ1tA3uTN1Zdny9FCYCcFIEOe+RgzXfF+V3rAEh+V3m2vI
Fx2lAxFiwW3Cmhw9vWLaifwTFdgxbip/7kfG6oypmB1HDxbALIHmgTweRXJ7wlmRctQvTXhPUvRq
dLnYYRcAXel8s642xNATa8RwFMBL3cNqIIVJzWka98MQjuYnvRYs7XNUaoM+TP9LLntJDGBoRO45
8di46ME6D58JBImSVqqQqbPBf5718uUVjx6U0fqG/bB0Q+YyuGj64Qu8ZPtN/YZjEUipM+AzwRfY
gy6so3kMtbjfL/s6KkO7X30LskbEMuPe78eevcBXiEyKzoBb2FciIy4QhbgWf6IXKr9rYLlzXpoN
TbCNJ8CpZSn8X+A0Fe2r0HiqcBDABfl2zD3p0/QwkakV6LrBvKh2Ml4kQ65TpbHBcnyBtUVLgMTg
q8upJqF4J3JfHLEFmWLWPIMbvHPv/H1GWuujp0qQe/20ceobxicZ+H+ympWH5LaYyuZVn1V6buMp
hcAI21q1BIZfSj+EIeaPfeN9aKYdy8KJchDq8KTYNFqUC8l0m0UR3NteSGk08iPI8+1LRDJII9kU
RT5AL74eVFtCYrJ6eh5nHSzYz6KyacopmDMfLXSelHTc8h7YaSpHNlcYsX1QUrnAFdl/cmrZV9kI
1ZoDzhbRuWorzhq2N/eW/Oz9TdEJKr2BZD7aCLiSZ/dA9p9FnQnF/q9vjdM9WXHrUKztGqZdX5OC
Y9BPOpJSQ9RB1/DbyANp4FOg/gMSJELrcBDUYKW2z/Bwhskv/bL3xCQI5g8x+sYlpcwAw3br98Aq
GvkAf15Z5G673nRvfvoms4dxq2mCjcrfq5UF1dbVKQnZkc/D3BiR3Dfw8aexUj4F9WqR/63LIhtX
G8kfr6m9c9hm6TJ2xlmEtSitQU4XL9lWaRjkjH+NG18mj5R53yW6BaKE56B4q3/KefS06egke1hn
QEiGKuuaHktvXhJt1lVOnr++CGaeK2XHyu7hnvXKDtJg1rxRof0A0JJJaaIf5nGAWgyM9x+sVNbS
OXTCacQMdNkqe9wIRRHffPGL+syxKO6d5lKqChcTDC7fl5533bDl+EBjRnYeKffEjr/9QH8rP6o+
r4KCuk0u3Jx1mYT8J5OI+Gft1qPYOkjJFZmhu6oywUw3TDazX1eFQzWRShnx4dEDFeNHl8NtXXB9
AgV+n/2Yp2KI99yq88EbrukWzq7WzYtnrjYYHzWjiCTpyUZj+oPvAs8+WmiVruR2FXreSy8q/HrZ
k76IuMd9AI3wzOZI63QtXlzfYKUjtXvIe7IWfJIfwkx0CFNB9IQEudSRMs1SVvybceJNfpW1d2LX
kKZ1/GFY8bSh3hBF9YEACiglqtUB63wemfk5RpWRDjpn1JopPQIgeJwnahTJb9M4lV0zYoYuFX6j
bBb06I/o/lkCrJ7cMDN7A5uH5qXsLkreV0KZ/WDiSnI5blZLiOa2wN1HDNtXX60DOG5vb061Bg97
aj6uM0NdKXyXWtt+WZcQ6qkClkE8Sy0sGo0rQ3rZLuUaFrfdGPVZbL3nkrpP4sSjAS1esGxJX+qM
iuZJJLlv4gjmp8ftPJ7S5bChOn+oaSfC67bMfLcKMbvyqePC1jNmr5ia7z9iHtqnSJocKLj8nY4n
bXaE3RokVT+mrYkCgDT8S8dDut7/Gj2ORv/tp+Tp80TyypMPyRHHJvMrXcxaWhmUQ/7X2spvNch9
X2U5hVwtZJYQut+5V7ZBaU1bhmshwgCBLaXY9GWuBFmOTyv+cEzN3XkYEsJojNLxaYrAa0KizdrP
SGo+ulzwgA61xxRSJ5YbFIUbPl1OUEsQtqTINes17QdfmqlH8QMxgBaFoGok1AR/19uOPqGaxD+z
nINvQVpTdxyno+zwjJmsMxWZEfLeyh5vyP7z8YrhG2V4OlEd6J+VFtwQn9jASbidFVLIzy1mtE/m
m99kCFKZPnxC9EbpIhJYqTTQXYrSo9cdBH6/bkHVlkYoB77s4d81AbmaVLdPUBut1RUwuut6v1fI
IKMkBGWzgBgMvVNa4JODtsjKSG+ILKNFioBjseDX5ufeOkThZXz6kIzdOCn6f7HkRhv3YvbtYq+w
TgwV2lbx+zPeGI67E04/TDaoVNMFDMttfHCeNgb+kSPQXC7LL2SJIKY5EoM24dgk6YlKmtm/1x8F
5Uds9NfRs9+kBR+sdFMUaCMNaf8v3QzvkbG6pC2MMqdXkIKsQBszXYfrX84BqaRsae6TBpRQs2iZ
buVHTHvJfyNjQmZ5IjK4fLV4Ka2qMnVP57SSW/QBGFNaSsmAox2nKwaPnSg5v/8736VfnYgN61uK
4PLul4bVYQ85Jkfu0qsL1Y/OCSpiXSNxdzceMeyVD2rV8DdYMrLchvvKSEF6wqm4TRKYXae9xYQR
ciIRVNzUGHgJuercne0Xay6A39R3HDWFz/tH2BOya8GOrGdmwbgfEJmoaVss7+pVTGFf5HvLSH1Q
IXOKzVcsjkXNjdJTdLHql2ipbFbfNnzi93Jxnf+iAGoAU8pyZc1bYFpyx5/GSPF1sG7w8kIgubdw
4gHw5XHQgJulC1APkA/tFVu79nFCMdOcR4eqlgnP7gc3PPQgtHB5eilCOKswM8QNocaQmglI6Hdz
ul/FRXwIdkN55YJd6mwUBbhhG2r3H0nju3tbHCczX7vtc5d6V/r4YnMwspJgU8h4YxdgAYu11v00
6d95hCyAFE7ahYqusgKtKRW6RUEE2sMxVlXsrUUYkRqGPNVxX58pwXH9rx2hyQanpS+6yRfhggt3
OAYD9zCCCM78wD55te21qBZgr4nKQQBSJeWFsu24JFZlBQhpYdGDDPh0CdDaWjd1Qve2nw1+yo0Z
2bIn4tk27Sx4eejcFluJ/QvRpPEsDRmOHc5AS6rzpiFRyeySCbkEGtATrsPLKWiOiQg9xZg1lNJS
WEw/jAk2pgZpuGEzC4r+c8GCK8Muq29/2rEWY69OM5iMu0RVat0XVa2SCHLvH4giGgMRgv7rqodI
Lib/5Tspze2Qx62sQFwDHbGMlyR4YA0ATe0fOxyE3LMk6M+4KzbSqWg8ey6qpzDX7e85rx8HZQi1
XUbum6RVS7NlIORP0/e53l5tPnayYyPh0a8r5mabyxqjby53EYxn8DLPtRTEy+ldBCtoyXJq3pts
xWOcesSoplahl3NHHk7JkUq1s0mmJ6jZi+/+xpKgjvxypczMPV0aol7LDcsRsqrJb7pZRsfpAy+0
BqM5y3rfGv9iwOKyVJQ/X1YODtJ/KbbIFd9Kkm7cHlCmCQTd1fkMSr43ouJBiwqhicKgxF+qiRz+
2sotlMu/eSuWU6cpcghk1FTiuLNUFdqhEKDAe3EdUQCPN63hJ46uPbumhpoyKyf04X8GnH1E26P2
DavcUPvm5XWQs1GNbjmJMqi7ONiJJCISbTv2UgmCJbvM38wWqkMAVYxvIoxbtyqRpzCgKVXL/EhY
t0JNWSxkCaK27zxZkFIwSKHPktYmBMMalzC2Cv4wcEwNvFwrzO+3wIetUTUf8A6kkuC01ZsD+fzW
5LQ2IvMHgYXYtv6hFqHhqnoJLW3m6bpkicl2e8Zjhwya9f5K1eJuq4p7m4wW9uuuByI9K3xy+EQb
3fuT9AfAJf7Gk8ui4n59mIVkQ8iLwe4k65e/y5WN2OGu8cvgSxbTGnfoZNpJqDQ4SV5WumRpmYUT
uSUAHr6OaGWI80MHxLd5WMc+jEifMTA3UqvcYPQGPe6uj6EWQP5BfrFeVKTi3eeUaniq1VqMhLcz
t5klUDBZqF0TPyfm25AO5onOjUltEzuBwLLjw5roGbFWUGc8IzEYDDK1QG/37G3P9Ns/Kvb6bl65
7iplDX1YON8RtUy1S1ay/+XzaRjgJKkYdGPRKOpTyhmb3Qzg3qwrno8fuRSLdvkDLCgIZEHZ3YUT
HQV8bhLWG8nZRidKs5Pvegoaf1O9Nn6KT4ghwAHCjocQudvzzGcMHnpslp/UyDXdo6l5i6nA8/qn
XHkNSem+PvyPE2Kr4e281R//Mfe0X6rm9u6vblYZ/YNFcrDdMx66AcvQbx1dcNmIA7CebrSEbzBx
nn5Fdqoi2cEVRJtwedbtMl0VvCuS0kDzG7unmKxT2fpt43KOx4hOg9palYHsxAlR64Wbl0qqi7sy
3tvdvRrJdchbBYJNEiAhAYqNNNF6l8NerDftLlS4bGEyR57IvBt6MbPDdO8vqWQGgDx72n7oEJUb
7YZcGIlvZ03gaNrV1drvwWdLFQ0zchobgw3uGMnZ5Nnr+HUlut6vI+ti/2bZp2w8aJxoOZ5AFVZd
srOXBiXdCk+M/j0/YrEI7eaxgk18T3Rk+yqeChCBccJV5OBDWsBqvx2Y/QDlgjrPoCFXwz/gsyJy
rqP2MF0JSJLkVtdl4cuga6Gh4vCTLfzn9J2kdO2ZKZhjNh2Gi1XX9WNI2xM+ULdY+4JN3zSQ0m9N
KHD8fpNnZXrYD11/9TZfv4BWztumGEti8b5Z1rw77tdBSpI/kV208t+2l95piLok0AjuXW4gfLTy
Ysyl3rQd8U6ZvkUYrbWoggWQa4dtvYvjsxynrAxMciiDUvlqIedHN1ucnPOyxVJPlIny3HQHs+H0
cHxQVElPWQJGGehYy9VwFTw3GFKKpGHzXw/W6MUos/iEK8QOoWX7LbgHyVRhSXvmRswezPkvrcd0
o7fuGkki7I9BqJEW6SbHVYijT4bec1Mse6se8DEFlETbfGEeg1TolrE0Wh6TSKCYvChqKBBKYhie
Da9XaoJE8+475q6fsYKPcoPmsHZQjLKq8dWavb5kHjxq4+TNo6Gh72fRPq3QwRHdt10sAmAGBl2s
mjejFr7eToGMjerdQ17RGOjRC7+YnMMXprXLHiih3LB2SZt88oPfXwb0hV22AhWUPDLgA41wPc/i
uMwUd/+JrYBNQeqSInOhF300VR2q2y5Z41C29KNOUF2mUki33Sysh9bH5dUGqJcTMG0PpSMf2nQd
QUidfTWWfjzwMRc0zn3fkD8BPxVFzAHfRpqTSM3IrwjDzYa+GFLVWVwVmi2Gm/PNHPG2DEUH7BeM
0ppzX7gHSnivYWva/WNj2Ar/CM6roGhITuJw+gl5bmB+i/OmWkoh9GFDkAB91Izwyz4iU21Wh8wc
IEk0AwFy1ILnpx2Olq2uyItDfDV+LSGe8EJ9dGvQoeM1/Io7zzgVeH1mj3SwWjrgVD4dhTlCGSwn
i6LKT+OGUIw8BFBkO/7MarerhrsELt5Hf2/Rua7shF0t5Vmn4Iomeo8ez+e1B+vZyOF4/8kex/6y
3THHaJ85TETOZAZgoTkxqbnXyjA+jM4S8JeF5/vdJYhiUhigImgE8UU7jpjOYwhXeMxxl0mD2jUG
3qrsfLRE/YVKnTj+dQOJObd3aABv/kGuIS9ZfYnLvdNWItistWht5G7832tcGnzXS3XYigaBD2gQ
9vIck37grOKOgC00AVexoYFcfiq/33kGV4hl1kQhFSxn2H0+98uZGAuQFIgYprUHzLqemlN0Ij5i
ewhIEcuyfmbvMBBN/ld0eOR0OFkotxPzZsf5PxNtAgu0PCpFfCmnNsH0f47lTA9bLfz9VTR14+td
kuM3qpen5JB2LAc7Zgr9v0xIASKY6YIcRGhFKCNeNHgq3rWJ7++1zH2Dkyt0V/6hjMuxFTs2EiZu
CC5TJ4DT1O4ihw/n4Dysbdi5TivecDOULmagWV8NDRIHBPbCdlukLcROmosiPUqdNN8OFjGRM78t
IkMLKSfeClV20VXUABT+Jmv5b9UitNzSzk9UHF/3I6pXEnFNy0psuR8h7bfZ1ctCkgpMaQm0c/sn
aEKaZuDELzMIB+C3cbuEr+CC9ki+Jt8dqYH/Hm5VPZ2xCMPW+10H+bttcUs6qRAeqkou/6fj+Dgk
vgsDJ5EMi0QwMRGnzkdlgutgx0PgVcuj+fj7IBPs/4HP4V93LwC2OuWpgbK70zkHJXihCoDtPTmg
IuSsKp/fbzMU0Mwbl7O3teNbWJpRzPloW6DGMjjTgBaCW9zGy7xpzGRQmd1s2JSF/9cWjVVopYfL
LlQKPwojWy5tioYqltDNrPvXmBHG8nU+ydYWpHueyYYGy+kdYdx/38GfL/ryx8w/rZMRU/g9clPX
DIQgVJesqei2xmvGC5RKcDPJ7zp97CF6R5BYAek5TDF/XXkI5BA/zECVN3UhulpHPuag5kVxdOU4
OhAvQH5Z8W/DT9vOT2Y2c2Yo9KAWxz7x7nWc3aI5vcm9RgRLAZRFh9US9sfO2GHdAACsg0ZLfquJ
Uh+dydLoY6u3+3orVbaWdS2DMVH3QbHDi0BN4xfvYmrSwC8Zg6dpUevBQP64SlV7GuOrANlbqbAJ
LryMLj8dKCdFumxLoGtUkvRKs5Py64lWoteZo+Sj3Os2fp1dOvGVZ2NazGMynJ2HmQjhuM+mcjYE
aXhqqoyuHSGv/gZ2nuxQa/nm4a7HsugHvM7WbH2sruTn6rFxWORLSP8O5YuH/5twBnp+dpQZIZiG
jIXqjZMZerhdiTdb987O+6K/TmZjGeEfSOXt1e1jN96ZoW5tZVMrteErwTVY1rgXCnsAYO86dGFu
XvJDpve+zFJl4rWTExzBYIrQeWaPf05M9p0c2nImWpTwRAzAU+aTr7ncMPh0/6H5b9fdJ74Udoma
QK/GJ65lkS9tZygKajUicLX2fvwB5encdSZ7KboDSrBfXZVXCivg2noOWtbZPyJ0py/RhPo/NkKs
a18PM5sX8dT40P7mXhuy7lqwwWc49tf32M9oX4PckXZZkXHsc/rT0Jef9khyknRCfH07XsxcUZCe
cRrTgubWhsErT7VgYoNDHH4D9VW6QF8UuhTbwaVW6oyfRKrfsecibaxdzhAXW4yhD+xo7QfOq486
aJEPEvZ0v3SpC8FIoMR3NKG23GUsLQ6wA2TSVdcgGZ/0PqNi37Ov7aHicb+ylV28bQIJynfcdVmw
M3vV9abQvhwoaQy1ciGqFqJ4JimSO7Vs2bQ+Jt0VgDB9eyXosf+xNbPIEUz0dTYeiuBAonvgRGpW
Gmt9zqAhpJW5EncyXFDkGDwnNcoeqitgbX7TnAWJbiIq61q8RCXjqNEPsWyevxvsax4wP8Ijams3
gdKR7gSyyUCqr3nBiw43/02u764GbVRlhyysv5LTV8GYhiBX/tMcstqj6IApFbe8tOxzFylnqxY7
q3kQTOH31GrUL6NfPjuFaGJSOzZuFbtQ4IG5B6Bid47KoQqGCDFnsAGEyVvXKbmca3R+TJh43Hkv
hi1PYZmg+LF456zai1UL6liBjB0uKt1zsy0ArXTRLUkxy56t+IFgYLf00NkbvEl49Gf7+KeYdgCf
rkDVQ+lffUOojo8rshD5fmKsJmL3UQcR5GKgSn4kNIIDHwGaaCn0U1mwuKKQkwp4qvJE0sJplEkx
SFZpm0GDS+SSq9lQL2Dj2E/WliNRHocPyvz+Icyy6VEeCLcI3eaXJytFzgqxMLAFz2+Eazs+Qp42
XA9AJRLQVNrmlwUmHrGlxXHvVWlH/XKN5hJ13iaBSVxai0xqBEpKc+1dr4e+eVTy6nXc4Hv3blPi
tsBhEsxGEIUE2sZd6aCi03GwE50gDEvC85aGMn3K6ex/bCA4GcaOy5UBHS0ZY5YGjEAZiY7oJ/sm
ylYr7R1kEi5Agy4zVsq9LsKi89PX0cWoIFAxP0pWs3f+5Sqf/7KYgLWPW3QHlTN0ZhRrezMbOb2s
i3ZtDoJfEJpzIAh+YUo3hVu5ojVN0I/E/XyDnMSIlJiiEiDBzD62oKeRZiQaebEqlIuS0br6gLDR
w3WTvg4LEbsIwWgmELoJYLOby07PwPgRy0T5JczGRlrTqAbpr5muEcWq4IrcnA1HOKrGd6noGIiI
H7vvI/IXdywLi9XsDrtLm6hup83G4180js9gdZzPJqb85JsIV2io0edpoyijsQAGN0W7ng89m2TY
4/uGL++VA1MzxvEMEuilo+4RTm2xo5MxwlF32qnOe4ki4ik1kzSBnP3tEE3tmqifsL0hFO9Pp7jW
3ec99gNPARb8C1MnUppxf966E7i79A4yWAtNPShBTi4H2BYFoLB0B01rt0teVykFu8Cuepocgmxs
fUpajI7gNrkbAMPSS+8SL7MMjwF72Rg9T5NzyM0JffUQJ6mXhpkF4XxNcKa7g5sylbGRSDV+9exZ
IqId4WlEsPTgoVULegQ3aZ3HXPWNJMqhUF/932C+33cGVSTqrqjDZVkeYaLCJbb2QzS3cSp7wuYQ
iyLgY0yWIiqruPWl3Ccuu4sXDJiVX7j5HTtyGtgtvVaurCvnAi8xL0F4q2RPaCRC3YITcNDHwDXu
P5fPlNlf+BJ7gNJiU3eu/8Elj+UjPbax97usurMvt1fmmkwtU5gEmklxzuKK5mPmiyL9JlBNqPPW
7rfCr/3g8jgBtNzp1nO9gzbbkQND6eTo1Ejtj7Ijd8C7dE9ysAlchPh7m5Rhda+Z5o/SaaIVMJZ/
ujCOcRLHJZsjEzpwOkxWTZQtIeJsrDS81tppY+oaKPwjbRzXXIMpqJcEE3ERrxwFQ4F5T1eC9wvt
zNs3ZkanMRUcO0jw/aROgGbnbZeH9pv4AQ1k9kTowgIScFkty4sH6vxJxZbJ1R+qXUT34caNrH68
XI77LKWK6Szyaf2zR/FiTBgYbgwmDjbM8VKWVuuSGc8L3UnYvlMRYVRRGjiXj2cVao3nxRcg/P3k
RHohNwAB72r8tjm+3ucdkOwRf2zpmxj2iJ8aj7pZBFHpuHSOfZrVzZ3yVcHoroG6vJDs3rnWn74z
kXitnKiKiJgPAJ0CS62Wj69oSegibPe+J4HEbfSrfyP5W4S8ouXD3dj4LEnUlzkSPgkii8I/9QT2
zhQxfnb/tZzgBztsTC/xXv0vwo1g+nRm65FgycdVancaXcahaNR1+6JO8UO6+GrmmMYRM3hQIdX3
9CnsWGQfHLy5ldQa5s1dqLJME4255m+Nq7TsUMV9OOecZm2WjVEW+/JW1TVxij8H0sAtVXxj+qGz
qq3FjnOCZ+crMkIm+xmCCw1wBGbCj5mLkyF//r0OkhpwfiIod7B1CE1nx91iCDsvWMW08uCw0gNP
8rYf1mjG95uQ/R0n4rXw4nt65UoClw4pHs+bm9M5wphHe2aGECHl9G+ZsjcrFvVWzQy2P24tnBYv
S9IyFRyprRAI6SVqy08ccnpp94NTJb8CsjbLXSdCLip1hpdQwouNHSGSV0f5tFwrQoazEyNtNhzP
zm6EBQFMloxVpVGf2EtE3XO1ptMQfIgnPEYB+2CL/Yzx/En5U3/adLustpA9ygjz3qRS1p3tYuik
jtQhx2ocUzc3FF17Me87RvkG+QUWrniCsSNCZLPOO/PGdcvjugZ1jJ0VPIpWIC3pWY3hCTaieCP+
0FR/AjOlZY/k6NdxRKXenuixztCOi+ffxVCEPjUFsptUfiCh3Kg4tv87fF75Morl8DxWCm9I9Gsq
cAEUThWcUrobdF9r7iExpdHbKlgM0FvSYDA4lYSNBcJkRBAlGmAqBtW+zsi7Vt+wyuyy3riZnsBD
nYv8+dMelKX7yu7rtNa4YBIi/BTV+xVn6cPl+gzMk0l4EBpwNaq9MuzMXujAxrMRv/pv+y+RDZiZ
ssWvYtk/baObCEgdwt/tbCi6KxVVpffbepjqyZEAex4IXn/1imwc8TyDQ0Lk/7puzDGU+Q47a4/Z
jU9AuHoeLQ52JR90PaAqlP/AlDq3YcEo7hcxv+SYne8H4+KIsl2HtwEkPr1vyXY7qC64YOJ5JG7I
QYGgvm3OSInzG8/ut/wyWaYyDgs/YVeCbkW51MXTTU4Yc7/QIOGu1024b7eufwY6cs9n6inOe9nH
+0pNyxuN5n3r913TlIYSWiAqUmbNQojhsHrqi4K2IZFa0chNU8yY1LRY0tcUEFT9Rdb66Wm6yM5d
xe/iS1qtEzuBZzd2ULlL3FnD0cybuF1TrHv9cJaEPhGIEkLyuLCiWISqYxcvaKp3EEUCMIQGyQ/Q
jO/cnvg5GXRUKfHaifsEEkwmhwEK68YyUZYoYozd5asxDdgRaCqs8wNNdPIUxGJu7UFQ0sXAzLjb
DW9CNxtAme/GAJ2+ccLsl+ToDaSo/uy4St/D7i0NWZNWzbsPmjhKA54B1ry4YGyLmT9gcMWwD3Ru
Pi7L2+mA84CVG4pkRwbeIp5qe9nFiW7v/PtNwQRbwni22XWnZ/6ZiPstnnwFmYHCSwttmGhE6BTb
6T4Jrqx5VZZlI28LktxBjDeT2M8BlgovWgViDLg323oc0+7ODVQ7SCC2fd7hhPj2Hu6slOf+Om5y
v44S3pk30vK8VtOw7xk5a+Oi0hS6LTcax36SwjsTchiWkkWCpCEJcfO/V/Fd0ZGCSSVlsirQ7+R2
Mo6D71tedI25dPKz/2iIzCdPrtrb7WcgB7VRQ+6nMRtiyAH2+S8lGFIiOEpDQGapLfADDm9T3PCH
EhGqrW66asWvuklXtkn/kqthLw7glOTnq5WDIONJN8u4L5uXOVE3otlXW0qzwEm0ux+QOVJtoKMx
1qqsAfQ3lvgvHd2Fn90jUGGJsh66oR+tfNSQNoGxcuGDlG5L/vjiEqZWbN4j2vtEVO5ouyv0YL0L
8SUKMB6jUt99X0bUR0q86EcCn4d387TaQOOzzrYsp4zVFMg8YGZHDyBr8fcv1a40sq4HJ6CG2OQl
4xN+yCdcdWmt8rE4A2647f8R1d/TKHHYg2RtmFzFruU3Zo/tFZqIeb68NXk6jDWqp5yPTb9YdZAJ
NCri3mpABbDvWOyNhHgPWhiKfwyi/BZiDTqsU8pswK9CzDBWK32SbnqNDu9dw5fwLYLvQPIoq4Ms
nrdxq6nQrJScIYjE6HiSg7ZQco8tuPX1kzHCCVoLQvMFGOxk+9Ih3Tw2elpDu2LUGm3zt7e3ny/2
EfXu9NCv8kq2pHCwH2s6y+1WkB+2eBig+68Qfday1Ll27VgfKSI1TnmCHfLHz5dLWQTZ80yAdY50
dEzVWiyJwyGlv+0XRXPV/4WA4bLmpkbWjXrmL7kD5OOW43FZjR1vPZ7lv3c83Jz0exhKVNKsHwTs
Ti7LmeVJ2ut2DKfm9tnGltSWt0yxyF34DQ8oUZCnqOiA/16rp9ibCKbAOx/c4u/lVAlpC2FxWTSA
Rwc8WFV4GAleCPJ+pNmSNOy34513QsLjp04NANtfjk8Xyy7YkQLcDsRb/ZQBvgeby8usGHCR5IFC
H/mIhJUsSU9JVKjWnVnWrfCU+HSTLI/obpQvn3No/Ds6siSjTe4D+HJZkcY6fVj63F+wUrPrxUjT
GlIfS4cpkTTS/EPcMsjijUDwo6KQxy+q2z5R70Igbl67Lyoqs5d1YJCB/uAGUwkNxaFKQYpajwKO
a1H8/BvaHwkST+/x7KfCS84va5CoZLb7vb3nZwV+xHnv/Q1MNmjxRLzC/av/p3kW2YSE1d08CFJ4
dmCc42q+rTCbeBUxVGUFaCkPrM3DUv2Zab/NOFk/Z4244HgWWA5MeRuSA1JlseM2FZrSfMzMAOgH
rdNLRUby1XTAmgOGjwOPT+/qHyWZGEn1krkknglWfP+792T5zzghbSzKQfPcR5UOhZF5r5F0B+7O
8GN3yvBRRJacFVVqK5ckeuNCDvpibUBAGrnfp/2JlvTro/s0Vf2XVnxf2t/PGwsNNaQ7rDyPgVkt
gMOFbakjHxIk8D0DK0SOdAkZBpVABvSkh7ujCcP4tYDSbWaI8o3FyRPz+nDbEHKxej4/5m6mDFZ6
yBS/hVnovCYEHOrJTHChrAHGYt0X3vcSxlumweDjaTtZw8jloipe2t7KZgAUJwnNZ372A0oRRgrP
/rkvwdULEPBXW/VpEBXHtYVEs2GhCz/j02rNxEQEqLnaTYA0SA7NgxmoX6J+VFU/uvCNbhrlkrfC
leblqlIFlHo3msXL9jKX8WEhW/Mb+hg4hcI1tT6WqM9RCkgZ9gwTB30K6NUpy7BkWUq4H7zXdMBI
sanYb/7/NeJWNq5k/SBtlhDxR4x5Xy24J/KhNoci9jjAOvnd9KTBqbO/zy0bVEkHMmDL3JhjNUsP
UuHBQmPue96vR4MhMKWkVL7v7cXDqUyUAYMmcwGY3Fs/fwyWEmqH2XLlc4Pdnrbk50PTVsLlDgmI
NY38xhIgdVV+1ebidbCHf+d37WswX/xT2EtpM02x9k2xIuSwXrxDEeprBUJXbw6qeGZkGX6wbFG8
6oSnS0Lu2swGJnUAtTkkMkg1HJNx4ZxbHtAb1Jdj8kD9NtDvBjwZXuuBy8y5lm5ABKM+xtmFD9Ay
DybPNA//gUlFcs2ZV8lYIQRqvRLlnY4Jl1znYE0QTpa7XN6dI0LygJFdxWYmWj/btaFC+BP+YJ8U
8Fup0i5ze0GFhS8atEvDVCuY7vFyN8KJg408trKCx3tCMejL7JMrsypncxaMz5H7Uza+g5QLhCvK
M1xjIXfrJk14+nENeIww6Erw3OAg5XQL34CQ7b1VsyILUzOtJzVZAkyhEyXl2QTV1JmUt7qg8KoE
ZhuLUkVNtTKQDKCmykZ6fY/65ymEq3ng15UcxJN3H4EGwJdHSWt7/KYoPUcZTT7UTyiHd9knvU44
a59El9Vj+iY71DTY9RGxExGC8x67KvlZxvTgGKSrWVS02B/llzYOpxzdL6y1o4WNUD41qoyATbgu
6M7IspaEUlaf5W4g5XU+Y/rGcyKHVgniD3W1dvzeOnpkK4XcoToprvednBIeNc9RiQF65oPcviob
T6DjKc03YLmSZL0N/cEKqSNr/MPRAQdP/QIZJbvskAMZezdzpkRRR1rNzvFbpib5zaiL7GkuJXzY
kuA1xUZArpOskxzhBDLsiAMwMEPU2v2b7NK7n6qoWxc7c04lraqvJlLqNNFbu6FkAbWFDaNz/arQ
rW7SvwdeL3qf9jB9YUDfJN84+RJS96SnaW5t6kkujN8e3Yp9VAEzF65nT0zlR4c3Zc0dsNrgcJkb
HABocxPxL6NsFXrvWI4qSdhkf41RhWhApMgXwJIntJeRKKKhhHM6KUpr6jdA/x7C/dkSuytPd2fA
n+KNHPet1no+sL1Dve4TAoKjqYzGtrTk7BF5G0rsc6b3rZhvY6S0qVs1hY8eS9bmbHYbVDVFABw9
rjlWqJt8atynOExKtR6aaokCw5Ib2FcYh/14Uv9QMJ+LCl6q2raApzp7kG99Mi0gXGUIZx/Ak1mx
DRe5kCPOKqs7NsK1fSBREKHIKlJeWQXMXrCrNxonxLD7JzhAq4z/G6xgLfl0QpXjJ8ey4V5pTkeQ
cEUvhVrZI/ivf1cSKtmwy8H3CfmBP1w2S40F8QAxqZyaGDug7W+PBrDpg2428Rsv/lO0+YzJexU3
v/k+Tr9ep7H01KM0+0cmIkAh6DuUnKdQpoP7YiUjYzZQ9ZUQI5NXr8a+XjLP/nr1Fn7fwxek/F37
uiiCGEqkHnSYQ4WGx31+gu8MOt9tp7BBtXmKaDKXsPQYUZ8SCyKiRand/awqb5wbC4inOiBGXk0t
0LGwveslMBu+jSIFjv757z4zhNV51Qb6p2lE1PTK94RkuM2xTU/ezG1OUMM8p/OP2eA8uD3Jsl0K
Rt5YplxykHV3WEah4kOVC7Pw/nyO/ImHKOXHpnw2h12ZIBNTcqUo2TyLNs2ozNwQ/GyIY7zTkYEH
89Z1hNfavYT4zqdMAs5bOe4NBKiOEVGK9nFmlHvR6KbLNru7klHr4Hh+Xc8DkH/8ECpvcr52qfUA
C66J737fKvz9fOuTyZzcA38M59Cw79XyTGaSre+ETy0jW8hJR/PQuQ/59kiwv7QXy8YiVg3+EMrn
sHNFPmKK9YLINveiTNAFsF8u61YlCnweokKkV+zv6AeUE35dGqFzFcIVw135+rik5rQ+z62jgEHm
xK6lc0Cf1f2udHDjhsc6+FTQy0wa/mPezfYBApJktg7nX8cax55jRvr+932wDZSgGEL3ZXCXH3+G
IUd2JfxlfSkIA5aladSppffERxk8ehndJs9k15+pASMIuoVwLe5JTYsjwTXJcdrDJ/a30ttqLmgB
ky4w+f41lCLmhhMEWFZJC5/ivEFJg1YOqmbGpMnOhU94NkJlW/34MdXwZTyamKE7Mj5j99iNHPmQ
kisnB9ZcRGY6BQNiby5mvpA1VEuk97UOKFt66bV/IIJ6HK9SeOhJJfl2Iqq82MQ3WHXLPGlObarS
DoBFtexF6w6kbsV1jz02WYg7fnMn8rCHDyEoPN7AGrd5KM+8LZiyTzOxDnXQy3ujCsQm0KuZS5zK
VCkqPXoQwEocq1M0/Duk3OR10CaWGqPfHOp9AILo+FDf7X528Eb3Z7nYKLiWsFjgxlMOLt/V4W2N
o0UoyltZWs7pDCnI1bRXjDT3MzXfmYwXtXnVwDiRbwHTUtbOvD6P+sc57JE8w2xvgLSRHe4H4d2C
5F7no5zTLHK3Zjqam1TUXiJTHYRIw8G0XWbUXc2INjoQktuDYfYeYOKR+g3yMLp82eONqtaXtCno
ghNbmrH4wai/Z1MEy7BVah6G/C5mEnP5+1JIvDTpVj9uQsEY7GRnMaMDwQQNqmin0mNRWry96+wZ
SeVEjlppYodApQczcqyGNZvB7ZwioV8oKsvSPb+Tsq9HZnp+SYqAO413jpLta62EAsilzhPrdUi+
FzQaxt4yognTKUQLpcCDcIYQIrpO4uTHiHCEQK82YWoNnDV50PYS0mB06ajYSzyckQebcj5kvF8A
+760eUH8LDA+r0zUhqmddI13NBlO+EbUO6SP/kFGtJ0SiOmXhc4g0l3xovOA0HXGrrcQB2x0XsT1
uEKb2lPh6XrHycoeY5P9YJlPfVfxqK78KYKtG6PtAj+aMpuFculWnMk7YWpI3IJK5yL+oHfEtIFZ
tpL+gmXISxzRWSa1doYMfhNjjPFSP6yl9nODVzhLg4XMUYuozRquqRiz1Z1Em3j5O0zD6lWSyuCf
6G3lC49FMF2CBswDw3q/JubE8FwYqWbPjTzMqi9kqdmxMsyNCt6mQjSwodxu/8hs27QH5eHvX+On
AXEV7rWXXyXDLzbi4Qd3xAs2rA1tfHhmhINVMM2Rc5Q5bD7vjusT5YUWvLZfsaNcOPGAguaJrOLV
V+iZqRulOWYLyXTXyWOunYzz9O4VYqZas13AdLBbFsPRErrEy6RoNlr8zw0nKKKtK1DAF7DkzxWj
uGL8cOBazbeLjnouzmBqk/EZTR6HWo7XL9Ax2hr11nPh0gt2EEa2by+PN6RhUQbza17O5mCNa45y
RaynsLXGkhIadRHEbiQFn5GRYwh1Qf1gH7tTf5WGQun6bneekuXJwU69xlV1WAKzt9ByK/mRwGqw
PRTGQh+ov39bR1mAXlGabN+QrKLJZwLlxtPx9DgnZv86SxD49h6X+T9hORNFfcP917PnhkGhrCTp
rQcZmQLyuy7l8Wu7vtsH0CBv90W0WClr/5Q1I1nlPemZAHRhEJWySUeo8VQ20nmqmLqkwlL9wKK9
g3Mqrrcg0KYbSvS/zBknCvfjCODfunZa/VOwnZpKiOblenylymO4c9lfEoLXnMAcycZHZu3bh7HM
JmqCCzrC8AwfOs/7CkXTpIOaJ69U9tidBi9rn8Vpp2SXRSNoyj8mTXHRvBI4f4+V/6Mygn7KIrHH
Jnz4EeUzBUmLohhW0dvsMPJx2gGkG30Ka5TYww4LivNWLeSE3tqX06FBykcvGuGuisHT0CcQDxXv
a9Vt0Xzpbp6PMTIHY+sOXIirxItbfJGM1jr4e7uWzYndURdgPVxDP2CDq+I2kq8voZWGPCO05M9r
t9vuJYeISye+7oCEQez0bd97LvzxxY4mR7B3wM086GLOsBBLMy4Va6BNXzjtQI9ZxMNYczj8RWWu
7q2YDe5oyxNpvGT971tlbKPaDSyDThGz2eW+vHnNCyX31dHfBZ1b6aYXOwLu0vNv5ekoIWN6KAsw
fPxOF0MabxO17d4GYu/ktU1zJEXTv2BdPD3vCorV1RBB5Ww6X0HlqLu3I6a+UwOEW5UehdBnXGPk
1lNADyMafwhYa0svVAyUU8NN+WnM0a/PC9GuuMYV42XeTca7SjjpVqkleyNf/h9LWWgextHAA6p2
oGzmlqXfYbBzAr2gKKIW+ZH0lrkC/mZW02/kKwmaGBf2p0SOP6sSzhgAB8XY2qa80z4QgcgPcA8Y
0KLNkR1cO0vhIXxvKyEsg3g4LRrq6ivK5bjkudVyzg4nGXU2jrkDRFr4YBp1C1E8FHImYuTVh24s
+brVei6FMRwNDkJBkQfuTdI4hlnFHYlPURPwGxvbhOhPp5L16n5L8kI1k/WlNZLyqL3OR93t/1kC
Uuw3QiTJWFcoBNVzrPp0fIbjTzdFmmAZCfLPYdOB1Z/cbZZeLZ086ef61ijBQ/Q5/cPO8PU6F/sP
Fq1op8Q81Nh5/+SYK0VkBLs6V5aaMmXdIkV6E4E9GtrB8hhqixdWcSt5HpoHqnS94h1Obd8UVNu2
ZS2O/jEDslnjmniEf7oGm19AQ3Q99VAc3PnkhwxEbWTTpyUfObSMYQLUCHKhuspzBYEc0zb3cL8Z
e29g77atQB4hJwGD3ldeUFLUiVeWQ3loUsbsRj4wZYyZadI5ZuxqG4XrDMRmfG+M35KR4YxWlZAI
QkFemqW2B82ON/TJ6yLShb05LsK6zYgMN0hTCVuE6jvpTTYF17NC4M3Gmy28n/QX+6pNzD+MBGvX
4d7OkFxvJl13SbvtPAN2qbpOzG8iscn50CW30nVwjkic0gDXvz+qaRA2QhIs59yba15jjM7U7W9u
0AdsddCkpifSx0Ixf36wqE0Uq3CwLJrO2YtOFUtn9SjLv7xBt7bXC/0gnhtWCA9hVW5a2Clr692N
OvgQRVPFW2ZnHArSu5eRMbjeB4kSo8BYr0JeTil3t1VnKKoEQ2+TUAizOZuc6ypMQzO9cn6DOIyW
G2A/tMNRHgHE6omwDINJ/ZiBKyQmvHp/f5GHHrpHlzagveUKI9Ry0af4GTPOHuBymHFkl4nwyThb
lhtXZvvPhWNBPSK34H58c9VE6kmpHQd/nF83Kj3bM23LEDrVyFKRW912MgfWJxPHOYg5svI+Ttbi
ulCS9T7j7n9lZREVE0fJ7evi+3mfthGDmYfa0P1UZTbFPg7CwgjRnAEtzwM67+GPp67KaJeffYCf
6yQqfjUTEg7km6pJUp4VPL0+iauv2g2PoU/4mhRI4IJCMufkp6jhpI3Uu6f6QeW5otgdGFZwkHnb
Rnpr2tY/ss/pz7uzS0o+nfp7vAdIDU9dy5w2pHaZpKQxrRbetKodBj+HWsNo8NhnqJm5uSq5slxu
cn1NY/46J7qrf121QDhkbefQhp+edNOvV8ymNVO+LL0tjokTUZKPzNZfLD9foPO7yKkObi7sJXiX
eZAjbGCt6JOwkp3QSaZy4xL8QTVxtjcSQROkJ98cVSIDKeRHYLaOKeuwl9QBHWmyVhGepeQyn1O4
Ic3SkFk8KHKi60DvXomuod9S0JdEKSKeKxxcYNL2mqHJd/bRxxZ6Qem1NT1LL4FoF3ZfHND1cz0f
i50uLlBg/9JveD7s9wlrXBWBTfYAuaJQEc9Hp921AWFMCJOCqtDrjPPM0blqxoulHB5DsTOt/tMA
3765Yule+pNYrX0c/XvHO6uqOCSqWMu95b/4TwCQBEx0UMX4AhbbdkE+VjswvSvD3I364b/I6XSW
R2Fh2CVJ1tlbJFLjmVyOU62IR1GcvWThHK2W8AiI/2TDweCzi0puhylna2x1oshCIIy3kB9uBj8r
3j5WhZxcaujCWN+JBoV8rK8JadS3RArBa/ib3XkD2i2MfwVeDB4/Zp3Ssy2Ic+9HX4LhCiLdTmHq
DckhiRPkiiTrJbf9BxTe8Ks17rJ6afiJrKLgZOijJ5QRKNITToOu6/0auqIvMjkBCNBYSYdP6pcD
RRyJLt52TVIM1Sk6/bsnVOUreeYyKimqV8DMuMEuwYJCI5Guii/Ox9jZ/Ciwdg2ouqzyVTqVNK4h
EKzVKbmO6NlfyvyHbKuVoyPjeItlwr/oE+i+PCN7+jpIm07n5pz6ZUPbkrBuqZ7OzB9NWIx+8EGT
rnpZZNLYouS9VAFmcHM+CjJ3rU23aScrzmkMlzVXDw5AbH8dRi8QHQjJcdJU5fpVYqW3Njwf2sl8
yBxffwUckdfQRe98sn9Ktbl75p0gBmpwf67jVnJp2rVYWHvKgOyqLrjIGFFgRI4lDeMHWwUY34h9
oZhdR9UVbLKhjWy2+7srFG9VlsQmpidCzVljqYp2NJN6IdsFj23iVq2At33D+Kl8cWujc1/WJo7A
ezIzXbe9+HwvtsCB10mgc0VuFgChOaspxZfYYmMXbgZbIsvN30jwwVx40UozJCrV4pNigogcLXQl
TsqG0DQrdYhOQnuvVKvvZfZIcEL3H8mgPFdKSgofCz293YdYMcqkJASkTKd0uJWfxQkQRNTWsXAd
AaDc9M/hyVkvkKuUqXeYKK2T45g7XAmrV0P9i9yzJmmzeBpW8QEU/iEjgmpmNanW4Z5wGFWO2932
++LnKiGUK5PkMfOb5byz/rzIEGWiHZb6J5iLv5oDO5BPiSdTi24WH21MCFIDHQh9ToXTRfi6KtNs
1R4lj/J1YHY2r0mP8Ni8VscOBwInuDNt8rRu/pVUVZaQ02xhduh8e4p0aUU0q/lfqGw9TnF4pSnd
shNialj1uroq9YGgrcnrGZZb4isRE31U7j17JWSl2N3XwbBjbAvokY4V1nsLrsH4TxyEdC72d98D
nn5y2g1pqHuUu5EW/DxksfRi7sPnlErOHms1PMAGaFZA5HaHXOxisQOf//nBfGnQyWt+tc/pifDX
1dlgj46ESMnMwnw9ok0bCL5tnoLYX+e2T4WC4NQsYXGp3Nr9kYYUzTYkDUkrObVpXN5nuYGxi0SA
HD0nAO0Zh3FQ8VEV/0XWGnePbL0+26Npzj1dBajFgzXZHwnTCuDVZIhRwadW4YH1ZZ9HVXRdGqro
+CIpdVjPAzwVy+AWBpQ9P/D5xryEWFeUzOwJISfXhG3cTGSUtFPG3d+mLT8dNNBvj0qYuS67rA35
WHn9B+ayVp1DlI5P9tZ55YO3EQcE79Ffouk7Y62Z4SGKyKQx2IHXopT8fSVrBe17TOAG6qC17h3d
epb/a+h0hA4GQ+k8zkoLluZdAnMRqsF6lWU6mTNIhuWC6WoTrPRAtFPIbZSWTr2xDlBqh3sY9l1a
ZrVWHgVuTPPaKur5qY7FW6OEgzBKLiZsBlCFjmY1unIAzrxwbABStRQYSZUmQEi27fQTrCneW8Si
nPVkJVwahIdf8hB5SqcR0PFd8hHwak9UdRy4iwv11CjStGFASocjxGO6WkVauQ+y1K3OpFcrJzSb
RdpC5m9JnWkz6xZsTU2faghbGriGNF37lI+mnkZ8hzuS/ronbKU4RIlLtAI/FqtS95GNvOUk55pX
krtglOht+OJEpsTW/+//IVXz8zmteV6dJuwr1KtOesY/XnfF7+SVYMTM8iDBmLaoQqffg5pY2eN4
KMkLdNIuc2TXY5zQBtlh1wj2fSZU0MSGygW7GNvAEfUJYYwK2D57ZhdVau2nBFOkx28rx18SB6x7
7dlTYxhQID8SigubwUicIsY3/UnGMuWdkuO/OUy+o5DPnhlvmkx/G8EL62pQuppHiuQNZkPCQrrS
1maVHjTjmAP52Nsf96TBOWTp9Kd3bhuvRrAfAkO8c0QeTn6qHUaw6WLdYfXixy24/Ns3Gjn4b+FW
KVGGlqm+/ozaFkZBYJ29CyP0xsXdctRvT6gOhmI5Xvoz1KO+W3Ro9R/OpYMxesbcF4JjksRedZCw
3IGlBbXhoGtfH0vt16xFNBz7ZuLF49o1pQNikjGIqD1SLzpR1GskhlEwGqENWBQBgyar7LCNOKuC
FkQjIV8ZHU1VLGAQVp/w7J+ePeD/u7z1NKJO/9xK6Fq8ep2kkr1aBY9vmFOaEix5NTLEZq1zn2oN
IngICaRmBsPZgBSldPbeZ7O4HBVvd6XrhY9po4+tz1Bhp42ohlJ775El4WqXzB7BgcyOCaY86O05
vj/W+fk5gIrllKBX6W37WU5YY+CIRr2OYd9hWGMYAP8dANYv1oNiUfxUjAXopN6FP0bNDGF00pM8
5ZMA4FE1QwCNOHOBcYwXxgX0FOZiXMT8hUhGFtUh/c6Jx5JdU6Xw02ital+hckrFUByg8iLgRBq/
f3LYs2DvpH3cw9jKHTWcUAXrTmMnGC7hmOMDGaa7zmeWnSZPq1KL6aZb6nmEWqu/PHPVWbrpeZnm
Y/KChj+iSwBtDYLkezrOtj0/7n3AsU/vxAuNsLV7VH4XvGo4ssoggebsxAnIKaHdNvjKNA1OAOeb
EbOcBQXDeND2j1Y4HL3BJ+FgZoDI2V++1JYCRGh6WdxRZGWZM9Hvf5YXCz2dPIby4Then0u48OOT
j+vrtAwwXZKBtNjIhKTH+et3VNBCyB/FNpMr415BHQZ6yhWBA9BrZL4eS3XrcPUm1AFKsF3WlRKJ
z5bmsz68Cgpkfte8HFiH0ZxgEt4CJpm5aXd3qVdUOoBJXkLfQjgS62myxTTvybjQhexsUmyK3DtP
9fOLc0gC/wRzln73MiOI44nfHonodDjC9GaeJOSZkKPAynNhqza+BPjq4CieZqEImMXN2jnMPYDo
oD72FtHx3T5o4pvUe5XuxtQR5L4uJ+ldl36TYqVNc1w3mj9POIATNkQ2onlNCB4LucZYRL8aGswp
VrwppjDUVJ/k2Deg6AVGNXvwEI4gl9WE1FheRdNGbu8i8M6IDXdZOTgFt7nKHGTBArHcf52ZAAok
wsoVE8xJIpeYV8QCXU/ucd3wOoUJX8lDM7Sd1xU9Wm/2XlCSvg8wt2WM2VHotNeaMt4SeDy97ikm
OLP9GWdqtmUOlkdKt/kdRaJeR/QpXCtsnVP+TaX3nkAKDmwiXLgzxsAi3ucUutjA9cHWPy83S29I
o+Yht+wAG85csyjPI67PXSp9avisjaw4Q0dRzszDAlURxCeK3znr4dAYIeL0rxsOAVJrViPbmNJh
4cfT6c+dPA6lTrT83yoXv8QbgvRCV9vEItRmm7DzTtwm/LfrstkaXGCu5f//PCqsfZUyj6AAznW2
beJbfoL+r/HgcsW83/vK/6pTfFw51HKthWOWVGZbAhOvhrZm+NxnmAGp3aAdCxWOfWvETXg6i2nk
kAZsmYVB9jKqQ4vOy9lItJ/xzUJi0rsdxJCiBj+B/1DMfqI/pQ1Hq++aEcIQrhxq+VEaFXPDi4/q
pi7ZZ7bfrR8L54ueF55XRp5MAAo+MrEhsiVa6rhuoLuIqq4exP7a6j9tFo3svOrwNlNjSojWM+ag
C41Gl7cL2bMLWrM/phvffMHfYv68id5u6INXLUQl1eFmQ73cqBjTpMaiG6UyalNiTYzoj9r6mksb
V81jSYsD/gex+bmxT4//O5+Am4apIreRys4SSMMxCWbsamJr8vy82pBccC+saQy93ZRrfg/X08/x
DMgAh9RzAq5eVECsw73W6kqskFRUC5qNFa2GsCPcDeUBFnUn9VPK/HFB4gULntugSA93VcVvd0ds
0FutUC6Bd5u6Aw31fC0S30n4ijpMSqF8fEVU8C4RzRC9GW9I5fQ9IouFxk6Xvatx4WIbGGz38RPu
H8hjcM+pFxQAKaDISFOOVjGZDMTWUORSO+ek6a2G+pDh9sJpIg9cJXWmiwfZ+HGFYPM1P+CQyy7g
qeQFtuRipjLHCH7YHhFfRQCUeI1bEKtbyWZa9JF7oPWSQLIDKWMYnD9PzkTXx82sjg+YAvyCL3Gy
YOMuPgOaJhwbBeMK2Ljv4sJSKZE/7bZUHD6qfE+WiUr3rKPc1ilv5LePMxmBXTwf08fuFxwzk9om
irgyZCCXINNO7rI/vZr7u/oSG/GS8KA9QySjhm6Xsuf4dhoG2oJFqrJhqhHyzIxFnXewCGDgHIZJ
udhHTYC3m3jG4ZMFLG9WkdfEQWTtdSyKJ8sc+Y4xQFvEh1JM0VoGXbHCwtgQXFjcyd0NMRQHEv8a
HepSpInIdzZnhgpIa341mJ3Q9+3xIJiezaCKjCrhUnnldFUU+qWWklCqf0Xq7bSPdOmqLwhpmG1r
5UlViZtgvwAGBkrSBXnm5Rncgn/44Fi9cc5z1Z+teIVo24bSHyCj6W0113vX0AYIlf/m2XK+QQrZ
gIIZmtdrIdi+DCp9AWvgGNcG1np5FVNEU3h6welNTStUDNvHSA6F4Lo3WhzCykqvlb1vASqL7k+m
YCdrlHAsTFqTXXVUH3TlN1b+FZZ0TnYqa5lVkSQPNO0YmkZTDf9qBqQHiJxMoFbrWMupYaKRsPlN
/kGAPI8Cff2kJL+Y9YJ3+nBQOteiG83Rac9Fk9aNOpcJjZa/Uq86votyhBjVtjD6c0zfPFhe0Vmt
6ezntsQBHTDH5vIZVJgL1OEvo4dkgXgzulx4/QUFBPN2VenrIMAn96eccUhk6a9mPTo5wQAJSsY0
Ee7ati0vnwaARJr8pTw6WuzHl2vnCIFyst2d9+UOSlLDoR7t+SI5T+eUSnahwGg6tObcTWwnOUBW
ggXgTmzTZ/lt5yVOZ/S3kQvDvgZN+Ca9cxeXKqti3Je9o1WK8C2L0DmKsIrnYhDc0XiOvxa/liBg
5zomY4j3RyzjZF+4zqubkZOVXyDT6ig7VhwGTfxDdzy0eKyN7FCY66I+SfHqgW0efMpg+fKlFnLF
oSSZCS5BKZxaROI7RA/5mXxgxnMdasnQpOFLr24/qE8mBl1/fnXrz1zP4Fn3Fw/rqEtkrGPtWq3j
hDwCHXnhXl3r1n0xGEvMe+OAnGpI7Lr+MJ0sWORgQ19s1+UuSYZGZZ+8/OfTinLT3NaHnWeiZv3S
00UnQmNADAWnasriroUJqqYzsj9gktb7nSZivF8rZjgPCSNP367U1JWKkXWBRVYSnSS/ldP8q8HA
hYxnEFW3b3vxXrV8qwPyZnG6QFCaaihCzrvII3Xtgng7tDkrpPe/KOAdnXzXvayXjMX4Q8kbIbHQ
+k5MjFwoGDWA1O3giEDUmmaBGofYv0gaItnmEsdq/+nhGJCz3VmLIEyOkzvA2qXGAv8BUipIvb3A
dwjFeEe+v4BapkPv1WWeE9HVrjw2wZjHMN23mk8aEarx/OQubiDx9ZE2YlnCXVOh7BBLGtwX4L4m
HLN4bfUut9YMAO34lTFw7a8sjl/3K24xrvUOrdYyRGYiWM50oILyENSrLzBimioY5jBrHLVNDdYF
XUlt/OAWvMaFVXOMLYexqmWPlddi4WssJOUB8pMTT85iKKtOYdFqR2K8Sz/A+YCrCMhea9uSfEII
9WeWwVWKZIqFyo+2484njM/3kYLXAhF23qJGqRRswOkRrw9oOqegDeyuGVNqFRWt43duoIT98hz8
wozGe7t46pTTLNHidwWEINN5zoHT2Oif7VCbqH89m18gnS3nLTSo2GQcC82SB1pvtC1gdnWcR9Pz
2pWjuCEVQeXBlX2MkaEs4N0w163Uapq0ZR+c9ntM25+taRTFbKrXghY6oWjoD7nncJdUjqkTf2HJ
Ew0wEYMuFe2ho6Sw0W1063c/LA9sGWgtqit4pl13KZXHilmRKWQVvjj5d9/r7cjGuUiVOPePIzui
2fGh/XHCfI1bsquE50AUU9ipwEjk0HbkDhYytjvqj4XSHwNK9LFDQ2KGlVW/Ocjc4p9tv4kcNz+L
jRjyAVUgaFkoNS3bfCsmn13L1+B4bYaXDlBh4nBIWFvJvPPKIuB2jjZNETozBFwUxQn26lrttLan
BLIyJvsm0Ub+2q9GVCSKfhJ5x8KAtMHVhPAokn4VmfC8P/K5QyXW/zXnq3yvjbNZ1OmaF/ifzgl8
zPMBk0QAjUGdaXn5wpjDpvzzAQ3Qxyv03ekKuLBD+0q5ZapoXc3i6zU7fUFFW9nRIf0iWS76epHF
aUr2ngkBzzigVASp18mneU+XK1mXc8PwLxPkfEDu8ax/rRE0L9nFV4zg/AdNoKlPLBDu2fRbxDCf
8CkQEMFsNcjwIFdyomaSIDLQlfUcG3pEtEoYzKWRLH4IR4bXnIaUk7Jat9N5Bp09LRx+q0AekIPx
ymArUpRLMk49N88jAeyBox/FLwLgZW7OHRKiptolocafj2TKzwOdW+OLOY09
`protect end_protected
