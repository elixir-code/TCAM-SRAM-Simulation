`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kOKe+xBTzF33257SHfV2ffZZr1PtLXjZ/uDy7zIT+hLx1+kMuM8L+eURot4ph+GlwCP0xnL7Qvk6
pLCEJ76maQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I7lWgddVDQVg9+uv3imer7WoL2JKEZi+J8SVKDYxLGYJ8n1E67ZNOeIV8KOog3gRLUQCQRVzQaIF
WabNhqKMnCZ/lHVlqitN7SgsjTYC1oIHorYaiZR9/hkSIEQVC1Y9jdoqdgL4T7FNVPFUiB2R5bof
vHmei1lsfWcDBK8kgXE=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bWFqDuIDTfr7UajYilTyOrmcrA0Z/c+7S9p+fCpxQ3mz4w+2fs7Vc/qHZHBKxBJjPvbLS+6Xq3+k
UhMF2mBNdh/TTmZ6ITTMZl+lpWkmHUtDYak7fbGHtqXd/SI0IVWQxT1+OnDypHRDzPm84mkDYjt3
lWYnKM373jFGp1dJUx0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ylM1uuxEs4Igzj79/chLzCXvbLbVsN5GccKhY2EYzWlwWYrRCJbxILFM3dR/SNKwMjUvUSJJcR5H
3vfRWuSQXZUvZGGiC3UxcuKfm2u+BdDtiXUjHnVXA61k52uq/FumOUHqnMhPmg1mQZBHo/cyS1aR
tw3eRj2av5DxOaaYJV2zHJu+9VAtL+C5+66Gr9WD4zHVuvkN+/j/VolBeAaWpRMux1hwXNt4AcDz
pALxHQOyl1HjQnqSojcDxAWetuMyjDNGv7r8kGsJyYMPz4C2KRUWCQAvGKwflt5dMyjc9Yh/x63f
pyuMZVcY17Ee3aSRvcb1NdtJG4Omf8ySs8yz1w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DrOzLqXJlu6GOjckvaCMbcE/h9c2UJLEp9E4I8f4catANtHMq4+8rT0n2XGL3f+xOQyzHYwAnQ/C
8b6yLYH34zQTrXqDJMGqLmHbPGLLi+9l/hJgKyM2wFGKkrArYIsOxbxUFOGiBqwyp4pA+u3x+BSN
zpHH8BAJFfRq8oiFh0GiP6gy0VgCSiWe7Zedquv/q9nqKSwnmPKVcZKb/ctnv6N8rjPzp+4CqLxr
FBQ7o3sQZUVKKKHiJayvpKaJv8HErWhc/Y5vNLyZBM2Pmmkf1hpTgrvZhBXvqPvRPnURsYtAZU8I
v42d8+fx6HqMjIR8oRP+i89emFOkXujCXn071g==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SiTfJDphV/Fy2H8vG0KSyIHqPS33epyZ9dTFanPWJ0rgi0lf4stv0J9W8mI/hMjDLKCwvqAwHEMz
mMnZ0D9GlMpRFnP6ixr4mSJWQW9NKyGaBcrcveoCT8mJUuguB//npSPyE1l4zIXyP/jUo2fQMpR9
lJoo9gVzCzlDNxjcIgbkYhEWKYneMEBNCVz6sFLNXMK14Pbp54TT8u7qLmusuBcuWYDnntCQlgrX
nAyuBiUD8wFvsnc8vedmG3sd1JhYAYC5ywWpQWaU99HwPpi3LpUYQtvmVUc41BPyYlSaTxPstGS/
u9Bfk4lxcYexPILzL/0Atx3FxgsZsZysst/UEA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 119040)
`protect data_block
4qVtsryvETEMrKi36xw5YbRAk2g/MBauPizZlI05IsFy69ruYmOy7eDgMsLHLrdXzNaLehxbJyZS
KIHAgCF2HwU3NFQsX8y0D5kYOFhK6EMx5ytcG9sQxp5seT6lFga5pEhzSnYqjq/vMyhBETYYu0Vv
aZhMOl4y3rTs4BZ4jwCdwKYvpuawmZg1yM4++eIhsYaJFEh75kAA8DpI7Oy9Lyzxum1cuSEGbNKD
6i+1BRgWOzVJTzL3QGOSASzgIEEZ/n5jm7ylc37Jn4tO4M6a0v9As5Jhqq3cQcAB1z5MoAwOufe6
OeeKMel9pteOtxplXyRCWaUcbMgkbagNUJfdDooXxv6xo5OyjXylIKksYB5lguJ/zVlVLU/7fzcY
HFFEqQMx2tEMLECGUqHMZRSJI2J/SyYjKdRcb0l+Z9C1AjH4XwPs8wnFbZgTtfGDy+z46vIwWSgU
NUZY9e+c5xwIgPRLAHRMxyN/hWcEGid1dMoD8R6dcKIqQhINcGhkhHRz7RSHzixRU2wF2bpqhbHC
Hty7ICko2bgDQ8PJljapZPCa6UT4IJHtvsptdJtktPeB/uWBZm5SI8QnMnVEXJkZsbojPBVQhiox
O1Wpr6YkOVYe1hjGXsrxa/sZi3Z8IQuilkTXIyPbdeZtequfz0pzIN4zDLlvQfeIcngSAQ3oEyfb
/decJuc02mMjJ6xtRu44GEt8KFMOVL3CKYSspI3I5+oGzdppoCK8BS2QHufcoEu4y1nu3dU4uWae
VzGZTVuU18+LV0DUaS6Gl08Kci4eL3JHOiM8Z/ErXabgEJQe1SiR4ehoNPOXJnPF1TF418rst3B/
02MsemISYrwREqYzFnXv+qmivOkDKsMHRjUgD7O+f3ys+rvpLNSj0HIFgfkSZH9hcVrXrM5YjcNe
3a7ahhqJ0YofyRwbdD8gc9T20rU+KNgbG4/vSZCHDiPkht6xLCAs3jKdUxNQdylMIuWCE2TVIuUP
1e3RAI3GTCw3KGjf9esoQv+rtNJ/yAP4ZXO01MPn25Cy8kdukB9LmxJM+HuXouFqdr1MGiTvVyF0
mr+57HfvtiZ4ByxXLuT8f6KFxHK2WHu/6Gieh6uybfiP7vbxGcDictVjKMgkbVe7p8+s4aiKPIIM
DQXGSdhus1AS9h707sZW+sBg3uOPX+/4VpKGEaH2gBIwY8hzyXm3V482Mvm/fGb/BLkupE+lM2n5
nRkjbJOx5wMbreQt0EykRDUvDPV+5lwcnKAFzF5SI0/xhuf2jt0+aEqUgeUbZ9iqTm1B+JvRoNze
+q1miFBIwWGsvE62XSM4GOvqG/Z8tiNHiP78G8v7TGIz0CFCIGyk/8xJxkml5SLbk+tuQLFe+Jac
0xfZ8oeLunhZkvkqgrkCc0qvNpvGtdfzIn0QDwzHXOfcCFqvcHUoSfaw1zRyrTxNlw2iDLURFxWg
lqWj530GHDzGQ/XvS3VE83vyAf5YpUh1X3dKq2bAoyu5VLrbjnfX9HnPR9ntQuf1HKuYCmkDDsSq
/WCnzoNHQ1Xo52L7RMCSkMUgc2R843aaHL+TA8eDTL55dcYZOAnM8RbPQrGpgL2d54eTcyF5JiDC
59qUXt+YDKLaIYTpPNiInJpvUSRBm6Fc4VbOBdBWsd4VNmteK5qQNbrrT+XSGdgaCqqDqi5HUd4t
kbqdL/AECund14ksIwJMefrUGSBWUfkhx4gll6ExQ3kb+hzIcmcwx9kNLry/v0lEPa1IebfQzc7w
inyx/qQ3ZI/7OdFFOEpdxdvSxk8kGfA7ZEKkEHz28a96nZBWC7HeObS0Gu1JaRnL+XcwIHfu3dJv
4NmfD80NXt/CRm8K/NiWaFJ1/esV/+xuOYgECgui9S0aG5sf5AgDVu3hBkzdvxLcjzSCbG4OwrIa
T5khrdZgD7nYvwnjGRfLgRTMoc/h82AUS89Mag2fqdO6z4A1amiecbXTEQ2ur9c5zeRX+vD2zHFP
TQ78cQq16E5OvhFgHd1S4o/VAfY4gsMDLrvkurf09VH6eARudHXZ8/+rpiN9VVbcRLpH7LKkYf8L
chxo4EbOPpwMoYWrBhThIRjZoBapz5o+sGLyOGtgW4+8Fhzm+T4GsckezB5IorMdUUvMPONXkpI2
dLwq+kQF5KypAWknBu+JrgQ+Aae9+dl5G1UArRXWdylIo3roNHYnVWFIg3HR2F09prHR8sBVu/OB
C6NeY27+FP5wAMe6MieO5MgTOq3CZf5zw5/cSSsbyFadNcrGnvdeW5J3Hc3Y1TYKV6coY4/4bU1c
omYIRwiF7ZnUX6uya2+cxHpE1wcLRTKddUXbMeSa735Le2qXtkllQSlXBPtJdr53uKusjl2TjSAk
2CKJXaps8+PPouk99J6LcVroiObMxVwbIbtjDAF/MDe3KyupSnA1qH+WV5QI6rKiIjGGd6qxBbId
L8/JixXIZ0H8yoi2TUs/OuHc+ussrtg7MsbPXbZESVGhGqpvrueG+khN7SKAMVPizz1NCJOTMJuP
+75tL1W7taN9JRWm/b5Ao0HhsyjwlE6LW2ZweMr3LQbkqA8clermt1QtiFgwtBSaeWsB7V7MDmZj
ABrSL/VlyAE/TlzrEokdhIZFEVSbckuiXrN1ktcTIDLNpH5GU+YAkFk/tddTksQCFQvlflCpH0Ij
PrB0SQCqbx0pqRz5/NOb6qqKGpp9/hUJLyCRcQWjmTpFEu4OspT6HvGp+WSlB/XsIsxl95XCdozH
EH1DkWLteF+Lksk1xZ3fdLub7OGLg5X2xKI60DN9dUwP0jyuRgTi0YGrVsYvYoypMNrV8rT89lyA
WhrJHQyVdQ2xXBvb5lUJw5kuYInQxwJ5DCjtlwFvg/xjguW0SEl8k46MUzPX5VYq0Y0mLERSLJAB
cde+Sz6hyTn1Q15ImvlkwO7LQ+0SALHKFgW78CW7WfNVRl47+snLKmC6COeyT6K+iMXiKQKZYpzS
al5iqDJ36h9fHyIwlUTfFjA9J7skrd1q9R+N+mQHcGnhaeTQkza+dcdR0Hz3UdgC3ftwL7EGf+Q/
4Vy8vrPHNaOD6iOpqP5lvZ0bVth15Y2tXEFCGYrpwBsHLxPqRtvMGYQm3SmqZAVoBp0JIBj+nr1d
Xa2TmFrf+QQs7MGhAJD/COi0uRjKWslWXIfpc3sGYkhe2RYYV751whBHpPKVCRlIx8mMNJauCh00
y3GS6ZbqEZFIb+4dpcXN5pHdp85B2RgBpTA4vQqIbb4fmBh/szXkGyNhuUhFjotyJ+wfYOK5x2e9
Dqx/ua4XXR0FO463Uvt7pG1zwzOPn5OJDvpAlrbECJPJSvW31d0Roc001eeINGWjmritNlNUPbvA
zX5Fto3K+4qc+UlorM7mMmYwv9HK1U+0EBxo/FBNoOFLmmOqTf6/VMrMFrpkzCuFCoGgFN70llc7
FeVj6q15vjhhuwu0Gp7GjTFZEC2CFNW3ukvDFfnD8q/2vpP8oFndZrAHA2k0onB1h1DZ7U3s84Zb
TkRh+zZyv4fhQebs1rBm/LR2Os+Gf1ljQ5Ow+46duECXBN4SWOoH7y0AA1wVLD2nVj8nxbdHgsWh
f5wAXzxc4FrLQNfpJK7H3ArEjXVtlEkBYhnqufLzBZhNISnInzsZesgML9Rbb7Yr3BkY7zD9SCCx
pgp6AVUyKcBABDsXnzy3Gxe+Aor+uSgroy8fgJNMPespGBai0XwGC9zVDYzh6R8IAca68K2c01L2
qbidL2Cc7+InipUOBF218NB2NT2wKh9kVhdC4hynKMulswff2fnbn7Xn4Ewh/vBe9ZPY5pMmLCrj
yA9Bx6H73J0sRzzpR2kc13r1SDHJJ4Qa7Auxk9yCS3dQLZANsecRRgKmdVbzs2xXOV+NzkhDZxcJ
oPv32GUCk145e12dgTa/4pad++DbG0L6cxGXDZM7UvKv/Fh0E4+glj2lgAQl6ullcZh0p1i5IxgH
kyPdHjVFm3Zim365JW6qojA0KCxFioiIwv4UvZZw9NElXCvie+zwpufIlGgw14Yfpfgt5iAtLJRe
CxtEh7MOr61P+SJ/5ArVqdMNagMw4SPNmcAWeGUGKhoc1nf7iI5sPl3Rx7aQVPc9ptvXxzhlrQpH
hBd6juPkrKV2jao/tx2wVjpq1+mP+cKvZ7B2jzIl39GExFYbIuoAlv0uvuBzg7vs4aaJP0DVsHdt
UcXgypjyJQHtcVRB6OB5II6hSN4XKRLNOa68Zy36rO0ctvQLuY7G33UNMllP6kCEJJh6bSvuAky7
tHo+OiYSe3Ld2iF4eirVYf9ERcGUB7yE9jTlFqCMvZ0c0uQLFNczkMmqbDARh/ynjXIe8tucUZH4
BOg2pqeDGwxVthHqmfXLWaz1TIud9YfgppUShx4VYd4yskAOL3gHU2mxP0BxuagCLDBNUfPjgYlV
arOUV1QLR6sYndAl8c+kV3cfLAKE/Pgos8D/o5EfML+TtI+Ecz21unxQa0s+DP4W9SscYm3PT8xD
D5+AuAckWPL/HSlmkIMwWKeL7/22/0BxAYoeuRypstOO2oPHQMj+vCkJm4zOqIvlhyS9gSPDxqSs
ExYqDcRc+2V/g//t1AYsu0/jj4EtSyrulbR9YKhvA/xSWRQXcOBpKY+ovKWRMGVF3izJOm+Vfv4q
yiila9vE3nq3fEOCxmWPK4DswhcJD7gVFsGqgZxX+y+vROnsXW7GJdQUOg+82hfASczxhNU+zLZo
Ys25IIssR7XOOuv7H47IFzIKlYby7zzWypPOZxJiYzWLHk3Hl+DJuqOEtaA4bH6L1Kx/ibFQmmej
PqZLGaauKYSeAUG6lPNqPu0vGU7WgZ5F1H97tBY3CMcNgtYvxV5gszju3FILef85fpiWZH6ZeKrK
/9lke6iRbCySblLeaUHn9RBzh8rlgjKgCeE3Xrgv5SuDhru5n+hd/WDGcAozJAVFCdCdiUCmXt7B
6eKUrYEOtTdLY/5Tl2R1B+M9H+h3t79WboaaOxmw+vBbjtur+E4tqO8cfvaR/OzAWXvetNLYI2UI
Tq2pE+nG9qpq52Dwj1F47IIyyRcSHRZovyDA86sQgoZLHBsY2EsqQmY2BDdr6WE/+sMVz1g1JzB8
hnZwLfZVNzRg9FqAWW5Dg4eRugTs6dDlu+dvSkv3hITZbyF5+9hf6b3KcmBiYQkg9CLGaZK1Q/oF
hshK0oQyA1o26JaW5UdikOFMicxLBjVnto8PQoR06b+i40IUz10gI9vaMaXFsohZdB0lHh03o8Yh
0lLtWbGq/bBYCLsjpdNQUadqZG0HzAL3AmO8q+bLu903PBkXEGs51SHr1lU6TiYrvlD2qqSYkT3b
WwckRxwhs4f8MgI2N6P1Kh018qcxOpGg/SOF5tfKj3E0Vot+QFhp9LvX4Ve9XrSJKktOOvl5hxXI
gnOBl26K8Wv2yrY3+1SuOu0+fa3Xbg+7jQ/RXf2Hc1HpEiootKyUROD/Prf/zq222SZ8hZyuOcan
XDjdZUiF9hWpmeRYADfBTNIi5HRTeqpEJz8SvSKEnSuFHxqSCNU8ZGjr9SX0uSvwJtcEPBQ26odQ
oNG94CLtRlIrbDAh4buDfghAorizrh7IAmomZ3g6rJGTS2IFsW3oE9xxRRWODU2EACB/1bBqQllY
cKs/7qx2Qpl86jMWPw8GfxbxaQ3tnXd16XcGKcJmJgLtmahu+2yfIjlNHcH/RuwuQ+dOExMHbjtW
Z6byv6bmA6r05SJGlJbYzK5PZlKWqL595ZkCSix7t2lQatkV9Zz/r+Ew5RB32POsJXzANEQysMTF
Ux8J8T8lTI7tPPbJA7jHmXD6etpTtIWxw9c+ocgIGhEpEPly8el2n6LspSQH8d/gwHO1e/bV2I7Q
Y7AeZUMqUZKGijBa80ND7ztYmE5YCr//FUbFxhmq1NCb8bTRjmFt5S9oQj232f50TAR2pwTx1jVY
Y+8ikgKtZphwXkgwf6y9vIF/ZspfPrs2fPEN7TnKs9wI9q7rWd29OL/i7RhMvRgAqOevp1w9396h
l9i6jziJTp5rugqD2lyk+4hRf8tzbXPSlTnMihj15wJXB2uY9+iJJNFpFOipyMKbEAnPFBFuGuza
3NF5K0XWW+P9XXeFb2rLWC3NOH9+zr5m97YdbHuglEaEbWo4qpJRaRIMd2pfytGnlyFQXzRMYAvu
4NdEbSjOtLLGu4fZmqe/SF/bJM5llvYXL/nyDtpADWtqAO+SQHBynNf9PPZJmJm91WPA/9IDtRub
LJFVTtmowqu7OzgWSLb5/X7GXBIHUpRWbkT1Z3Bj8IQ8v+R1Z20eZt40iATF6oOk1KopMLQP3fBp
7dbguA76BA3oNBuqjeDdkP2S9dKZVZTKOpIUymaxS9/Hlskr6tW5whTby0E1ociG+BNMTS0vmgKc
cnGe6yGsv7AZ+Gp39WJ8z9kLbwXhq9Fnj8RlxKwQfyheZ7EC562Jm2fr8Ba9rn/mv5AEI8nMRV+A
mkfrV5sZHZorZoVcvigEjTJeZP828Nnv+xu+mkgWd00IKjkdH1eaf3Jx5/hjiORNlhMHUTc+K9Sl
r5adtQUAmPc8p3g8UyR+Rfi7QGLGgeoXHKrT1XE72oLQdGKrkl4QO2E0Jm7nESZ/rY3RRq0h85JM
vfU9XRO13I2BQFjW/zPORQ/Ne7eZJ+K/3utqpj0THjEgHuD1c7ZFwYPndLlEnC251W7Yq27R2eGk
WFxrkFbKseQKypQUKyCOa2SCFf2e98vVIne1Bp+P/xI76Gs3tYtm5JSsrK8HIhzAmxsr0zSZlufQ
b9d75995ps67khftHeTg9jWzd713E4wvOd2TQ+jaMW0osomuoNOS8HUvBEkkjo6t3UIcGtXNLgRV
NmS/jdRiwtN6avmvovKqMERWAI9mWRfj8t1Z0fqqdp2A7CLB8FcZo4Ltz2kvMwfF/+hfkmJV/JR7
k0gOPkqYoN21jLvXseGAKih7tL45V9nOYGxNDzMoWB6HBL7TESRmlRvZbb2uUlk2A1Gaw/0h/kXt
cpn1JDWG/TFEEe5sx84sk9udg6vQGfWsG/UUiHg2L764TIPHGxS7lC+hfUws8fnl8VXRfoPT0PbP
otj2xyDV1YjK3K+jzHxSgLJF+BKvHp0dclExc2yXOdFufZX8+mErOz3ajT0IiJXfL15t9J77VNYs
EvI03CkFWOLvag4h0rlkJp9pm3kMn/C5w6H7dH5GhhBNt7/zsbRl2RBL21zGosRCRYsP5FozJZSw
en1NaCnHQIgFlSwK063ozumxDUvkIRsT5Z2gw+jTf+s+zF9sHStz5CQjcLpUBNh5ebkN7dX/qrX6
46vjscMK11vl3Ha5tvJFkeIzdS8URneubPhfizqWlMmyhfro/frTQ6d/Rjg+hgzjR6sWx3fzob8+
9YTLFp0tva9Jh0cRD2lsXpxms+TjV8pQVRei0FQwnbeTRITarSVmJDTY0eUcFRNw0JSaIrzzMj6f
R/eEJ8Ji5Z6v1h8/SS0fyq/GyEZjkxVrJa5TK2km+s6GQ04GYOMlNSCsy4YbfeVvVZt9kpIFduvU
yBdWvI+XNTPJnfwWS1DnVIghRhD9arlSIZDIJSNOQGMpX2F7sYYfs2fU17ae1fxr/B0tyUMFwj3P
P9/0DDS8nITgXZXHYMc0/Wj2f+W/IcphYSPGtyfi7y43cnJaHZ/uZ2KH4gzpDzRgucquPdjXxlVn
iazJ6REBL1LBxj5Wb2jVwS/MVr2matJYSOyt/hm3UuZuZkkkHhtS8ErsnY3jdSCc6Eo/2pbyayfy
3vWA4PIsJkCAyMdckbjWJYwMAORMNCVNQ/E2/wquKvaJWw9UQ6rJX0RRGjYS+LD/B1NRcIDeh8+/
QfXuzJiNqi5DcYleC1HYrxXasekidcCv5CBlf8Of3Mft88ymqGscDO6kICS+7Ft0UHUDvh8VFsDu
3Oj+WK5m65luuRGN3Fn+Hq7Aj0UPJw79tgImHG6raxNHADHG+ppX8eZuI9VsjosA3puRjKjjj2+W
boC5iIF7kc/NOkwmWmofNiqe8FYOKSiBwr6nqIlMn4T8Ed0DHlH7xE0kMUuyyuvK7/AfNfAUZArS
geg4btBhAbDjVbUscEyM0z+qF9vXhrj/Xaf5KiSI3k/V/ii8HdS7royoWpPCnVi+9UK5PCJOBQK9
0kJihcL2UF5SgdQaRARgmAu5cUFcTd0oAKlBVR4ymuRdR88GzXzqapC0HAhQsGg0oPzCq4F64OjP
1dEr0ysr8uxl8q69FBROPVqtU1Xwc9CnzZKPEKdL7cjVC38HCZEfTrJciojMbMl7da0E4Hliju0j
Oin1hKXcgZxM5Do3RaCZlt2bdmglm71q8aZBwzzyjOSjATQ2u2xv1bnPgOcaKNui1K+lsy+AxC8+
gSZFPUpAH7Mh29aqu4et96hzT90YI65DnEIzsU0cfCz7balxzqDg8oNupf6LQirV4EJ98cu4xULp
l+tptCkmDup+LFQWHm5XaWCTGHUw6CPApnt1aCB+CR99Eak3uWIpznuIgPWwzBzydvsXNiz6fT5x
HWGSYJ5uVmby1yr7rnyg77YMRG8NSxDoHDKFXNIkty3jbiZn3X1ohbJP7coquHGYMYQNsxVZ2oBO
+38v49RG7zNMJ9JoOS83o26bGZSFY3Rho4zXKHfM7g+xzRHD5nQcDIBSutMYk7jMnvvdBcgC0BDP
gWQFpgECpDQjGvIlzKX9j7wMKV7eX/cyVveKRu/PLRgYSpz53LFvqd/53bDylduvND5SdwyjeRXy
T+qYyTRocOVGmu+mysS44QWlEUcCQscR4nMxXwYG1Oqcz6vEZ/o8gu2qW6xBVGT22MqTSv8bLGpp
qx48TNPgv29otg1YHDuL6Zbh/X0H2n/Krd3hcu0T78SXc5ETgTPf9cEBj/AfpRwKB5wW5SQ9RDro
vmmKg5skTa9KCTykiis6BGQjLAKYWijOgpHnbH0IlBXzULQR8RlZ+WttceDHezUMkmdOBsEKCaBN
W7lz3lXIe7E24WpBeoIOt/ZP6XrZHMb/m0OKLu6/fiOMR98JXyv2fZdsBnFtD9mr+Ykpk2fyuTxc
UP2jQ90Wj6Yb0WWLOxzCV0QVRqdKJSPesRPq3qA6GdbtXXRXjsvAooIPcq4NFdM1RV3bi9SyzL/T
ohzpf7OOjyFoINOpkOUXapCsvxneibzc6xjRHRHjTw55X4KZXhnjNTPxuU037M1reWzJ/2cMjK5O
8QyYsjd5Y3HzBILEz7sJcXAOVjxslbK8fS5tx2HIl0zjggHOyjhfT5Qu3OawyGZ3Ok512NU2jlnT
/imjxolqHpRcigt1VXGfCNfvP+qfnArQDhDrLIVTP8Cn+5wET5q1BIOz4eJEBsfaiVASYvahaGTY
O5lJ00QOyBVd5OEaxjka9zelf2KCcjEafMS3+s0WWd8uEkIdoBbc6BqToNg0Wrp9Adaq2Ccj3T2M
1DkbtM+u3DWgUKVqnQQDSUV/qxbEJ2ObM9u2g4JcauSSju5OBId3uUpq9SUcpnypknCJuIDEOSSf
Kn/TRPYlUT+R7dS6nEqcUezkuSISUOc5WatvZQNBxEyvbOFoV7Bd0LIHfZvyA4eX4B5ptoM5Ye3P
G7OWzDiXRV3vGPtmNaDq7FKM5lw6d2QahFIeuDzwQGZR9748tYLQMx19k5jbPJ4pl4enLMwxbG7E
KtEhUze5tMwpK5FQLgLFTEiOES0yBfMo0SrWPDGWdml20OAjJWr2yfVBJABnwizi9IMgVMuyy1WO
O4DPVQccoSWy6jI1+UWi+PbeMK+T1YkVCN10/wOsAvgdFqpidi5rfH/vq4Mf0Jhvk6OmgBncZfPU
QpmlA72lQLvCA2Y/Z30AHEIFFIv6Ysh+TA1ac1yPnoy907CLvumZO9cbL43KunsS/ihfFhDVcU1K
6eh+fcFpgYO7ODA0taZ6KchaEtCaPdu/7OMIfiHXfdShart9hp04n1yBVn1kx5kDK36dmf/dR1NM
VRKyx3iRBVD09mg2QKs4Boxkf3YZVDA6rQWu3YiqL22IB0M96f+3Vzpng+SYIhZ+M1Q4lGB9S9pp
5tBnzppA+cIklr0jNpWkAaFsftiK3Q+keF4V4PM3v+p3wDct07eem+MUpjfKJk3wO8KTgiUj85JY
bDdqsdu8Hg/Ebt17gRQo4nbZnYJ5CyiDv1zGFbYmZtwvsd9Bd8SmTjWWDW5azdUVMx6tyAEpNk1A
OxmJYJFuP3POHRjopOvq3Z3FK8Y/eCoQKDAw+6XdSYnsnbU6OECyeydCEXydU5bYkkc4v2AwW+uZ
R/Cx9ZnS+j0zLXDrDXUtgX/N/t0axC0l4qhyU/dOu8eJYcQUby386DhK0VRarbkcXu/8I6dHZqSu
LFdaDBpqaHBeQE0G8B7goZDkvaLPARTBUJCeF5ZGE7d3Ot2/qsKjRZaiIZgywML4j4EmFU5Wxccb
U+zv/gvYOM3kDTIalot6h2+AFS24lJdadF3JZ+C3LH/tAUGlntyXTRXqKFhw8uS/jsrmC74o75BN
+4VKHTB1WUG7dm5kSh7kRCf/kUWWanMDRl408SfLEV8bY8sD0G7JcMVk6dWxvRctod0oS88aw6RQ
/56B8mqXaPQ8HCyVLzN++tbz7vty7ckFFc4zPr5dRtZ7d4VQK2Z+krHy50NUG9a4z/KxIUCGZT2q
VjibCFYmHoKgBkQCsafrd0ttTZ9NyNT9WGwTQJ1a5Vqbavc3ifoDjlBquBOucZdC5kkNvxKy9dHz
b6XJddkSZ58TbMkcPKCVgRsCxyDKXjfqOGlg9FDfpi/JKGfPpnj4u0nvTy0kANmai0g72JMdwb8H
j8jCM0+A8iQgE8NvurrMYdC7LOtOI6FPn4f+hld/yK8lA/scpoAJc4XrnKU4mwOlltr5xsjgKmPm
x0wdk1UgYmVNdVlnewxpFSDBV5a3J+cSl6zA8nL9T0mpceCFzPzo2KjVKYYtEZgWOo3QiOfCAJWH
feTWYA7M3Fi8HBnBPt+ii3u9OdwTiWss19ap7ikzu9+sy+BxzImopEfnXOB3Ey+H7LWZ4pI4BG2y
smWXgZD+iurDDHaPCwzAWtj0DOBi4QZS9u1jaMP7AfP01pgbhNLvA9vdJjvPMYEkwriUPa+AqBn/
Vxrd6L4UFc7Q3lPSx8cmsxcbApuEFSKjbzB+bxCgG+UHdyA+Gzf/r+l7YpUMUL9C4fhyw9RFJ2Kw
orBdPDEdl6l9zJWHlGdeBJDDA2rX4E9rC6l1nxE7nO/klXuB1MEiQikqWijZkWsCQmFDEGiDq6mu
z99rDhoNA/UIjXI4K8NPTv/0ROsTdY9qoGyM91q9xEexrjTKUdiTglwyzHoZ2cFck7MEL9qtXqBR
gPRUqjegdoqXeAgUvAU0+cysXZrWkHW8PHmhk2rWgIRYsEB/VZhKz/A2EYtZokyngxWt7aJo3sGP
ZtX/an5N/0hWOAAklx7QGI4pRkYtwIMNS1Q5xRE8KPlsurXZECHdnvuH/ClJF9DCo933Ja2u53no
TlI3rJf1Xt09N/Oe1+zKvUyDcJYJ8/uv2Fxjg0AMHdcMz/asht1NM19kxjJ4/w6YEHE+7N2ugv0v
pbBaZZ4SvXQPgG0a1gXW5aLknsogBhBzzo0eCssF87BzfntBjL/Et8XUtTSeSeFHWy0XE5OUrHww
VngxvdJ0MY/mzAYClhqJpnsMB58VFmAOVzQAYwdDP2tBbOdmhnTLLgIiOJrXDRfi8gB8kSN6LSBk
aI+/VhKAQLdKGRu8I1hmqfr9xjdkUHTpKyDGBDbRoKLFgjKg8iEGth6Kri2VKSxMpzoPi4+shRIz
rYpIcyPIcvniHiArGNoNKH01AJcYvUwGtfkroLvW/F6HJbnPap+9qPClCqDJD44DUl/Cag3GQSI0
S3o2wE0laSt9fAV+ezysfah+uqNaQFVQLdVZkCwot2P9UnSAG296ItNX6aWl9J0VS7Po8bsZnQuW
HJviPsgUG+iPuQidsUrR45giL0vQqTfrOBLJSqSqLH0zncA0qJzc22rRC6dYSQkQ8y4iDixfvt+A
/QmGDyght6Xmq0kcLqwcGRqU2LAi+lT6kJyKg2oY24kOixzy0lDF5/lJM10o7nJzyhogVOw8EOzg
yv8d2PaYL4hZTC0vxWfPIrbuZ0UG0KGKnIXymi02JuRF+Z4g589mil5xxnwDCT/PFOCqEcvtXxuL
sVTAaPNfZN7iTGnr1RSkVh/iWeGYMabTWTLXNFfXLXQKgkVY3DPukxrPL4kxeMf0+r2jHkYnlaQp
7EjU0IRizvvSruoFmBu/vj0O/iqmhNhe3zlD48tq2F2EcB4AvS9Ze/ez+kjTwL1NTvFFnzPqD0Vy
S2DOF8sDfgaAr2r7sKtQ5mQFI9ixa3OUGJnjjsl/H21UIskmDrKLz/KgsluNO9eAnjZKc1SyTHNq
07eN6nK9cCML496QAHfCwWHadbbrhgR74qonuXffLdKJ/YQPWrxvWU0W21tNCwULJC6dNCReYLYI
PsF/ogxt6YWJJQ6gssbyIWTAn70mIcgDpESC1FWJq4C0sHNNlpo3iuWAGFuNIJHq9RkrSL2o5fjn
FnfI81eikcPbtqbEIyBFU4uk7XxDRH8QF+MaNoCvbaU8ri7xdhR1cYmrlRktywmVUbrVx1euOHbl
cbG5smEjRo3Tabu9ocMvsaV3WCgiefyEHnvHwfYStjT4QhorP6e6pBS5ajX6AVrYT3qpLXPGy1Ag
bfw+NxiM8jBJSpvxCU3NB4MNlI+zoQlNYl9VTRECOrlAsRMI9Q97cht65BoZ55msc6k2x+WF6Vmj
PwU+jM1jv2js8bm14nd7o3agKL1lNAM2ovkobszstfl70ckDv8Y6jRLUIareNKrHs0zY1K94Au+3
QcexKyJ/ydi8BRgntDlhnTb5jae6JJqfm4lWr0BcDeXBnSxWHmYtv9UpMaduU7RYy4enar66srZv
I35MitGBnDgQwvn4NaBLkoljdiheVO+s5FJgRVo7MsN80OKLuohG2ZgE2fBIbQLWLWvFTNtV/NGE
jwWOI93GQI+DVn+VQlgnIQVtZo0KBq4NgT6CAbSisxoJTUXnbHhVnKOrBDlAeRASmCcvYqSBTZko
OwUy6iIvzEexED5/ZQdF6B8WgePnUGpL07HrhAyIuAfPi8BIXHAuADAwnRPP9pwdZIFHngf0vjm8
X5DDZ7ew3SP1iQ/Ug/tkZvBrOqZjJUBZ8OOhh+Qlv5g7/TwrJvCXy+yqNrWDqto1GWV70IgA48Fr
QoCZbzWzTvTaN3UiR7TP3dSoROAH0J4eAxi8gwHTdSkAReR3YosMcGEubeUHzdWWrQGO83K3vAN0
Y77PsofbuQQhn0R5CtJBPQ5Y6rWnAq55sKYWupALjojN1I7MWuWodz3bkPwpFwfNZuWc//lQ373G
z12iD0D1zdiQRy1W4zXrorkxkRVQBhzAFuNmONKjOXunsC79GZ8ErqesBAKwVsfLQxXJYYqI7K0S
TThFcShdsn4Us5sQ+a213mEqPy+nPR6+lO7PKJlq8zjy56n3muMd5f3b4QUz4ivmmSuEJo3+7Dc8
/99ORvHtxA1veNJl+uBPnnOMXeLXhWM5ZIREc1N92MLDsp3Qb5uUa9TjsCZe9jD0JgFJp5JZnO81
yZQtaI5MK7Vr41I1qDMfprwapYe4zxzdYSNrYmFQe/Ua84usKeriihImJvqTvMyve0ZJu/cg9N9I
f20SIJ5wFDydZxaECeECuRkmY+e1NjgpWi1Wh0VFkdruIWWLDtK/o1lYqlct9LvIL8ndjTPoAKjY
EkoOjjvvp+7srJq/8A+9tqJJCY5fNUF9FxPaOoH6tL9vL4tBWoKt6Kco5jjZdw5EyNJOF7cxNbAb
fr6ThfLq4PwduhxwCVDF9Fcs0xMUNL5NYJgaqcBL4XQ/uZJWC3X5P1EYL/9ANWCjYe8TrDwT7hqo
m8zH3ZB9T8ku/zW8UJtDfoMwoUERe2v4PjTnxKGJXm9iBZB70MLkrHY8wVCxZQvfhttpG8fT16fm
JZjIu6xfZcp5FsxPrE37eUg7K/BCbTXQo6p6Awf+LgCAtx8GHWnCNUIA/o3wiSKK5luUiFV6n4qh
DOMhhgdMs5p6I1xoq6sP5BJ46z0LfbegwxIxw4IWb9K+THLV+MxG18GXWqFC7bFFy0LyqCgOn43x
XCBjH/iAL5adoDSlo03rH2aIpoJ3wcsRSveoKRMIhPLN9bp0tyvUfaNHCEjo97TED9GWXS+9BMuW
cnmosBjLYRawBV/GdtcauX2jnJPpPrXNYgJbcpRKZkiFb9Bd0TQtsHJaqkQrwYoaC432hV03/kEG
4sh1m9VUkdjV/yoNsXMyVuLnQer+bC9oddotIyF3vGLv1MkdRzVPpH3ub63NfZtMeako94xvE4qK
6YNNa+ugvTu+7Obvq6pY8zImGyHe8Doah5iCfcK99120wxIb1nAabZ0zjHG5upZ+jcr5P7SrL9i+
mtoQPKEgHzPFjsY+KvIffz1n8Dz1bQGzp9MGYqXRUu8uJAlJAryF0rE1WD/iV7XfnblevwOZJnRA
zhPa94J/QpYirHk7QS9avkVFWOfJ20FQqTnvTWQLPJhkKapHNpLbLKbve5UTIJHiqMFFsxHfSTxA
GpYSvA+9zO2IkgOFwt0F2Q4fDuiDV+pImZ1i3i4VHXM3WVwt9hSHaZT8bxmOWre1fJQrEDSUBUmH
MJG6xwIUFUeV1tzXS5WY1AphEOyXMp2wnQkFk7+Pic15eEsgBDjeb0RHMnozimqtNzjU2BLDBe7c
XUlSZkVyEWgvoa7FgI0RN58/O5svE3av7ODA4ihmLGkvLFzt3GRWSvs3F90NIfLaU8Ux/mlIGF4t
jVffBZlaP9ILYJDuHl2+F0wMT0UaYxwEAB2gykbI724UzKz77iNPP4IJO6Ll5c6TduVT9YogEgtQ
LXXxhYE7cLYjOYuF4aujM5ySh3pmuY9Hk8WjiOi4H4D5VnhUBO3AKN1CBlX1Fk5l1qvaDWEINzta
sBPAL/o0EnRMcoG30So8GTEb87q77TMzkzVwLkULFxaVKGoJC8mfyFPIXZ/V/BBlZlUq+oAUALvb
qE8iFYJynevs+VixzG++WBApA4vTo4oOxeILW4XMIl2fqUKdr/wHgzrW9BlViAkOB8E4otWQF2Ny
VpNlOkq2mDoMEpweWJBLSe4OvjaitzIWDL360wZ7Mdnclh7/bFPHR3rJgbB/RNXz18UORlTYBZBc
rZrQEWZ/P/JQqlA/X+jKKsCeAqKqZSnEiC4nD240rI7iJ4Co7CQ5pAdw68+d15ti4FuAOUFgNEmD
fHBeWxH8enYazeIw+w8Rav9r/nueQeGXj9p8dtMOhkLdjTk7T6XGOcCROJVmJWtR4fmNbVhYiqx6
uAv7lQuT4NHG9Pu5Y0gyly9eJrQbCGcFJikodRw7zmTF1TzXLvUfgpVSMappwty0kNzv1d1yalT+
SDq5gYycDUGFvy9LxZyLP33ZHJEqV+A6T/RnjeMkbsr9Vl5+9KYOvPYBwFnmNlnWnUOpnqlkhYC0
fKhDQNxqI8Cnx6IK1gpZbT2q7dlVSNYFaSF7pfeA6qNJGSQhH3a5xoNaQmWkgnS/nJH7zHh6Jlip
WZIf81U+GESoc7Yut4FA1FSuHMN5b2/QF7UWTK5i2ZBvK1d5ClQFKvJ0OmPwf3uQLs7IziXRXf5n
QnfD3pPvW6pLyQmR07cWfawR6nXKkYH+LjZDWf7ZFVeaXoHfVblBnFWSBYL58hPrSBv8kpl+dW85
DOCieZWjXOHMJC/KA2+JlNE+Co8oF/XJ9PtIwiC1OJoxNaSwvhkBn2lIvMt716qXb3/wK0gHD0mu
uVggXoHvM1xOcuhP6Qs+B62YlExx4fHr9unB34hDPE6he6QJTSQfj67uj+hdJ73WvvOsa4NnIZI7
k078bx4b3iUsjWbh0wmugcO8SwsT0X812+bpApkoKTRRQX79E0tnOboOONU4oPaGl2BuNhYPhKHM
uoSw39Dfm9KE4hZ8qE0EZb5nH6En0skH4wKpQnPK3PpO1a28KTO2cGdp/OauCElMTKt4JiLqsL3C
lIBGKT9qNHREE0Nlh7CqnMuTWhB0p7Juc211BETgwQlCGygNQMgFxIgFa/QiwGtDPaBmM0bUVZb3
xWDz7jXMc8MEbrwJsIwzSEBvPP5C7Ejoa4YEoZqa3QbD/3O7MyHPw6t0ih+qXpstDjkGw+d7QxQl
KKebdpi0o9Mi6Ro8VtLSH5HP9XXA8pO9SrHZJ9/UTCr/lAhMweONbOh3vSRJ6iMzReFVac96rjeC
hyc16RG7ai1bj9CtyE0z61Wu/sQAfPuCgiEpUUhVwWuBjPf0s0hQYGZ5mmIvT/7LwcidwVHNzxsC
KdbSlXTicJoxD4+zBLUuod/+dLsCjvGpfHuHNB8JLMOG2/lstXPNZknXBzHA/7cnzcMIAthS6zQn
06HoIgtuE0yaaRGFHalMYbaWNrwQX5MRugUtJEe0JPLgxcmeIv07Cpej9hy0SOd7d+GqyaWu7y1Z
Xguiv3kwuixRj7jGlajiuiOzPoYF0BJ6PB/Cu9tymDlA6oatFWFNoPf1LeOTqSpz9/HmhxQ9Sq2Q
Sng8rSheKJ2t2DWqs1rNnFGtcLXVapyHioRKLPfhdbQ0l4RUQgoPqDPceOTeK4y90s/BpR/fVQ3B
dzMQA0JF53Jsb5bGmCF+bSfsJ9ZgfyErYonT8wjDo9AMOaQVlssJySPUq5BtQk5mV66s8PpTcIcJ
LvhY5tWFdRghFa/jZWpKLJOI8/AgiQ0Iq/QFFs+c/YzDV2muO46120GJPW0rKJAQL25TYGVxkdsA
1msfVA4Q6zqfEmrQ9gKC8TLFppbgprLmFMMvyi3NvJPTzOx1+IYC7lTGCA9p05/W56fBMz9A2ChW
kTSGHna8K4HZT0UoNODOBo/COtIh/q8wMwemHuP/7GkBny7ZR/eNhWXJoZVe3mHFaDHNFTtz5gOb
TUU6GP4UgRiCS3l3H2k/oyoGPalP1CMJAgwCreaHOPc8iTRueNTGiTs96RkcgOJiRgwZZEJOQBpv
JnWNCnMMkcGpXnHvUEYyLcVNjWrR2HaMt3p5lNOL6IH0zmNzpAmuyfrW2p2GR/186gH4q6Z9mCf4
fKkQEyhSA5M9Fwi1koXOGVW4evZF1MEZWahxT3eICAhrS6uZp/dSwaqY92EcsP4aQ0tirSCnBe7R
oSqHmPmVeyg4rxzUcqngxDKIPpZV05EjG4vd5uZFCDcZSNfyt+kcFoMBJt0hI9kHNKM5kRmmciz8
tqIZ3ZwINcd9gCxOYxI6wsZyrzbIfP1SdTNI31IdyIVt9PWBetQYN0d/GlsQPaNhbA6EKsovaYwV
C6LWidBY5udefihEuP4Q2H2c4YnlV0bdasChXJg3MvlGvsifCgKatf+wp+esylyfgUiXerUl/S8z
D7Vd+TugEPDRz9uBRcthSVdQUL6OXv3x19Z6wicpaGVupsaRpqzFBz2eXdJUakFhDSYc51IJmlGp
tUBknygyZ3/ZKxgIBgD5nSBbM/ADBtre4e17wj0LD2Y6AYFcrROCjKlepiq50xADxBpYGjh19/qo
8aJ6ESrDS/UOF8Ira/WGisSOQ6s4VKGIHaDN1cWim6nJzEa96fJ3g8g4z2JvBTTd2TSEchrJ/G70
R4lVEQs3goxetwXOdvhVRgGIUMt0cvnEzj6Y5DE1fnUSWCgPqDmygXDQHGCVeWVIvtwyDZyArJ/B
93ZEvkC8wdZnq3/dpQzVZQmoSjf0KHSA3JBI7sN8ZurM2Aj5/pIxnXELX0kAEfXV3kfFKZiMRxpD
BNcq5fm2jMto+ynIhnbvqvcitABMoYx8w/U00velOD9rXiQjhHOaD5f1jN7B/vZa7D2f7YuwO53y
gBWQKwdtIBbMvOBZZJ7+tXU46Dg5KPC2hOekyvB1fSA9naiRbSX28AfY1W+f+Ui83NxOhd1sRthO
kTLxgZXiSgyk+QRBexOfQfl0aOmvt3DAZ3wjW4aWlXhbm8Bgbnr5aFTA2yiccdAWbXUS2f89njTc
8JbVD/nSIvFCbetBQoh/tVIEejUJ/uUG1JqgsGhsvj9JX6Q6AJWrw+pSV8J07Zvkh2IWAM1zYlJE
VO9kKc6COkV5v0a2m77Tcpju8P1U+3ZlMjk/PPmWJXjlP87qyWNwIV0TJxqzCgbQINxuHD3oyDWz
YCUx2hjhb7qqdBsrV1EvaJ2vPqw/NW6xh4eQbNVNh8gCuUlfMgNbkDxOuxuUZW9ZODx6cSBCrfnB
mFF053OhLYk6rmMLfZVvUjKpMRtItwK5lS7iPZBbbj2lIiABYSGK1Hl4JfFD9nXNzMK8PwbEG6ki
k8Kfax789Vzha21PBKVNhQK5fMbmJk7BeRYGPfyo9ykuj8A7qJAwF5WUktMGbvn3jdCzlH6B0dbI
2EJqStGgUMsHzvOCyzXKjnyGKwGq+VLvD6qv/PoeD1AnnuYkr9beuuuV6fA/euhwbhs9MgB/lR5F
aspBefT0ulHcmJEujseSBARwRh7VSPTrZhPuB+VBZYXJBceEI7gZlTbbFj9Vs05q++8hwiOo6bui
C+PBBEi1HEHtwCUCC/4QNnfwitfQVlVzs3bJQN0w3/UtvFk0OGxCwdds07pO9ro7i09DSgDmut9t
2lk/GN7DE4tvab3yNRed1JVF26X4DkCJez1k8FSOH6i+d4bJzt2jHEHKSSQmmAde75y0Z8RlwIk0
H79tAd5D2SIJxd6O0n69vU822cRi38HjK8p+CJtcKSWwDEV2XNmFECcu1EXU5J+KMO3ZzEmIdTdx
hFO9tkvMdi7fyM6Lev8QJ5IXePg1QPlJxZVXWuhK2pXNKB26LZkk+7gu41stzcN5QqszBYJnnnyP
kwz2nXiMUg4lHMV2aoVGlZa9mejfkazqwUuPhPh8X4oUvcwUA2BZJ1DD35NBlXhUX7Tj/P/jP7Ah
TQM+gQ9A8rZSqbVBeAOE1V1Sk1s1KGpp48qhpBj58cnOy7Pxz1PJ9ioXlGg2CDmrS6ArSNW79yMY
BhWMYEfJiPNlWRXwZWUiL8GMX1bGz/5XigeTVafQi1NYYuk4XBn45Z6tvFJXB9pMXQKmeFyVEHUJ
6yp8u5DDG9T2dG+igrn7xqF9H0+Hyz930o3BBQ0/BlpgEvLWAihj/ddUzGS9eYgoosbhrJZVXXXN
Aqsad/V8Mltw936RXaKDyCDhvKVAP2sQFj6f2Xh9FWkq12PXJvGs2GhpL2SX6ph+s2MyKuRZtBB2
zhTr3GiFU6ltFTc1PqtrO1BvIhESy3o5xuHbGFOIQb3804zqKhnXQaDugt3LYTkzu3JMy29ciKsN
mODIsvuE5Vsnpu0vmR4yiBrKGMlTueNZBu4xC1LkEVixW+7DLeORbHwUUbq7wfr1IGiKE9kXvELy
g/xbu2dtv+Fz9ftXsgD32SmL0qdBKJtJTVHbwNHhCHtGlBfX6IL/Y7MiHXlDVwIk/L2WnNZLsJpf
vXxzx0dKRTcgoa9ZacwL6LGwnhGd/M4SvCGpMgiPDtwDHl7Q2R/EkziMUV+WVNbsPXWSmr0Dcr83
sL6Z2SznrR20d5e1k67tVKo4ilnTNPjyfuE5kmxf1y0oVrgPt3FUF+9jVhF6vbYd1RyQFARojjL6
cu4FRsP9q3sTarc/WN9/+fJSvkvDaydRxNzUwVeFGaddP2319yY0EFhwYdCq6lDhKQv4k9gQSN1+
bRi4yHS5WOGD2yfiW09Si93uA9n37WMkdLI4S+G8MxDP3iv0redB8UjPXl1FSmXMa+tDcasOt7Or
vRKT2jjewJfpwzLVQOVvj+51t9wgNy6YUMBPb4pJawig1Jk20YgJBrUuITLVTESlsk+oRtyZxRa0
VbcJe0kIkn6L0Vw8u3iwp6bQYZgfeYzPg/5cS+9S5pNWIwEGMj8UbxtJwPFQq9Vi91RmmWwLOlEK
Gfm7rV6seVSln2Gb0fghQKXEHAncumBFFRxAi8IjNZdHbNJSj7H6JuETa3bMKBi65p/sB7KRcwhO
sQu2YBTsIgh6/JhvNSwFA1Yr8CYjOQ0z5MtnOcZbHpIm+ewv9Hwc66po35sBucKmWrUtbawCUo4X
8UX3TNTFYP6Ez3mh2bN1UGo7c2IsSheAkVgrVCZGdsoBBWcw+gs/nwWA1B/HrVamNwV0Hf2WNsCu
zcesaQ5CQcg/vEWOpU2Z4ORU7C10XxZoUgvbAL4snvt1XmTCVQ7UglEOscTrXvvak0s5CBzVgSEW
yoiyAFk7Dt/nzbqfXQa2z9+Iuz7TsSX6Iqb/pwMg9lPxk/ElO5k5u4LPrA8fTeln6xm+zvdtFlaG
/Qaoudfv+TLGo7zwTemVKj5MmhqDI5+9uCbwTgRV4NKGjwvTf842rV9sw2FeKbufj60hmM1uLfcg
jtO0oWeeTvMPIVcWlsz0WdTcE9mbsXXiGbHw8Uj6oL0LzfuEzSDkHCTUj89ZgqDLEgzwrB5ByGlR
UYtsQqruKzcnAbi5rpmtiIBdHYnAOk4UpMbKEZvtOIWNWVosOYc7p4gJD8Gv4gl3PMFNI1nkOxIM
8V8E1xekl5az6os3Ayc+34Oe0fnX+O/0f0xEeqZW7wN4lWDVpfNDhSc2FxriidnwJ4yfFAxDQC9f
5vh6tok9m568RPJ2vtSjlFMBhFhGNqyoc0k6I33OQLIYOhcumSPFQYajvBaFETB9IRgHI29HJYsk
aAMbPfGNKeACgBkRL6gTQXKFsiuHC7kKLgOBRa8vWY2BME7xTd9KLh1JriQWj8hxWTGqiB5jX/GS
rJBCP893UKUdxsESNKLp2YIGBslYZe8+ptiaz9Jx+O3r/fg4ZPacK5Gv4I4+c00nEaPYPDSxIi8/
6X/QGE3JWZQsgOOJB4y+ywPgx+h1m6m46RwUEQXFRVM+lWXZyZcGkuLTfquQDFtwyC2SxgMgDVkH
jJthpn1qkN76rk4lUXc9aroyxSNSwUYpMTy48u/qKROA9ZxQaFbXFWp0uXGsSMkpuM2nfQWXlmJ8
dnh4RT8fYl+23rQCXuMinEdJb3CdIqBh5g77Uequ+t/zyXOzEjzvBqJnVaDq1XLgVx+kY/CkwRh5
9uCTuBQ4Qo8IN8I6G9KFdzRqVFo8XwgSZDl5oxKHhT5E2pJ9HKZ5ZuNB1C7Xb3xExbNCn+o5lKND
0W6yCU9t9IF1hKhNtqtgkgiMTgy1vKTLhVtiwVeYKm5b67rpFt4kaTVvm5Vey2LCMpQVS65dpuJu
eNlT+vXxQBRgOqmWivVBN8qfd9hT72cUwC8x3O/esgbSoMKRtNfciMeQycUA1mvHMpk3tFAkM6sn
/QBSI2lGbNbLIeTQ56ZXbmIo/Bj3r6cqNo137/gfFLQwWHXkY5NjnYnSyIJViWG8NnIerHBG/Qdh
O2K/oboUPjhC+ttoK9oJsJ/4Eyz9PowkHRtXDwmaAbH/88jFdB6q5FJV9YDc+GYLyij6Emm5LnWW
VLoEhtGZpL3nVojPWzwGEMs2ihfosr80zplsLEz7IYmhcwg7Bhb5/H8GKxClrHKMvIC4mwXJV5/t
elAI/EAcVpcnXWZ63SswUbBjaoJlVqgpWwHVqmLGYp2FOHf8zD6UCHsrXb+dtIlak0KTCtXdOFlF
APjZYMsJXZLLvmqkLiOou/3hfcl8bv3Pc02w3yy+GVIO+ypBSKWrHRw9gwKTcATbh+3KISph9qVV
hzNROVO3bpQpiTHlgEFX49bYsxxpBCCbsQFo6bOMlfCkKCuj2zy+wFJHIwXg/bdLosq67vYpeEx7
3UJBYVmltfXBljI7Cwcii2dWOVcneKiEfRNErEfRC2WavdZ0bI4/3JMupGxomwaNaTEwa5Ty3Gly
t6Hzlf6MKv1MzoAI1V3LK59M59GhkZN4U2oO5AiXe9Bk4dlNHwrbb5xeYoZ2/Cg9v8xpoN/Zldp1
GR+c7ufiVvhHZQ/BChez2bP65dBDwQAZ17JoJJJuSW6DSdiO+nbjSOyRpihu32FyOVNdBBXfI+pU
/0EqyAyKt01Ka0UJSTE++iYTiGZyaoL/U1BEQ7HCr28LcaKyexl/wEwWTeu4g43nC6LdffWrofle
DPMy+l8lv8FOS0hPP0EXKMiJKhEFAW7cgERyRVtsN7spX+ng3Ym2P55bLrCvXv/1lllkZumo7Oru
iDHtUX0ULk7qyXyDsEnhrwJB+5zhDtgiIg3wniecBShg+0+oGTirQ2ZO8RqwsaJy62cPbz00i0az
q4pxtoviYlVR4BV7SncHaCQ1Uyaj7I7yW17TlgRH9cbDONwIgi1SQ8gTz7wRvt47AkpBhc+ObGkE
9IjbErtpt3J9Zf8wg0B34GfEiw26aLmu88gOZtH1fm987zUEhtQCRwGkIcgp4JKizybKZHJZM9Rr
uWnAxiyvVPMVSdCNfF7kIx0Cj+TbBuF/XoCsPBeKs9TUekAGEbCOy1qqMtpsiMk/2jUftTG3cyWS
cIMtLgQ9TQl7rETGjRkOCCZvAeLB4BRwibFC1aGTvO2gVlAFdplA27W77RBQPhqeqxyHBeczpJ67
FfRrpemiB5yPmuyQSSUTVrztOq3CcjBNPWfD2mfbzKfpkkb89/HKWRPcVh03sm+otUUjyn02QOSU
6/IqMaC3XWrx4O5V6hJ45BzOVBP0vzN46n08r0C+JTymk5AUmg3+b8bqCJx/O9al0GjN9z70nJaU
ouh4wHNemcw4AOMbZJxUQQ/SICxHw7aKtqxvHfEU493A/jctoJPkMJOBUGbEQPM2CnwhcSDqAkJP
LD8Qae57Pgmq5eUQRBdOmf/ITj8qM9thQWqKQKOxxsxiXP6mfz4UTo5+0aWD/OEpFJGws0JTp4Y0
WJVhLkQA4MfdbstGl1MH3dJF0eBEC6RRshOLWP7Z8zKUP2q4rhug/KeQYD2ShWICrDqG4LebGeGJ
mrRZpPCoW1OKN5uU1MsZtUDCPqHMeP5S3LU3GqMFkUL+Vkrl6mIC8BKDslynvY//3ooClPvE4kPs
C7GHiYM8NNj03g3mPkIlitgkk3EjnnVGAHopOb/xm3G+WhMIziCOgIwC4DojH2i/4xHenjdyrUj1
rkZ3iKsXQIVK7zzmtMJ70MbrSD69KHaG7GiAj5scsj630QX+ZKwN9FzuzfGCNUMw78fO+8ZmNapo
X2TDhZszGoa3WTjhOdORqN3U9YT21heGNtKbi9qihXSlQr1DRgYHu9s/3KY4pZ09az4jIsz6Upas
ZVG5SUJzNBvQZI2ttHETJgb4SEbOtV3z3at8hrh4ncASoYPGsRh/H+LlAX+qxyX16iKa58Vn+HhG
p6F7OfHEcK31PAKUNgQVOVjl36pslcc8sXBngUXbvy72O6I2Da42Ej/ubaDFb4H0eb0pZBgLcp5e
Y2Jua+peEKg6GSUyJyeMqJ85gT/3vMacI6h+sfhq/mTFp1r63w+w99iXnXzG4ywyID+orxVVmsxu
hNyuKscH/Uc40n7D/bllbpXqBwTu4NPgRgmGvZJ/+XPhb3rlMeI/7UqGJLHBRA/8UoWIYtZswi4w
uu9uECQ+LjB2Qp+Dj2ax8zg1FhYv5qJw8EHSkR2g53YlntE+lm6fsNSTrEOU+MGD5YxH/5fISphi
67bCyt8NKbK1UGQO5B8wWWccN5mhbiEFWoYgRz8BGwekxH3u6B7Cn2Ll5LVm+66gEtEvYyV/wf2a
3UKI/238UQgQLCKidyzeykOfYz9eDQvPguwpRwQ2EiZq9sJdNQIAr9kryt9Rz/HaVweOYRtDHmN9
ONMiJLpRrXmpbUMzjGdF81YdTUV/9bd/EFLgtsBnmfwR9FKCq2McxmIOdX9AWxUS73Tu7hsChh3v
Rnky8QHavHCM5S42IUYV1/0xrye6g245GfW6HBaWiHqQjE+GKZ9Mm80Yz/aGqMVekA1CiMKetP3h
IKf/WycNRNqzM1nDW0sEeG1KioZ5wG+DYmQXxImp3yzwKU8neZp7Nn7AcDoVVafUzwLIhSgG2Q/3
aNChvLx9JjurV/9h1P1pjLD721kjqahKGeM++IoS+j+H1aLh26g0kpnSCZwlu7CmuJmJZjhGjzl6
aNVCJmGIMxEp9laQB0oTtcNdTR2hPYLTTkYpo84H69TKItLYpyxrtrHdHB8EAe4x+G7U4wscWaiA
jnxHAjhsHXv5u8Q84rqnuVQXpBqipYW+CnhPp146SQwlcJ9kQWqgETVPyGAzurCi4DkYgC3lB4V1
D2xbvUd8+1b7J6qyoJR6qD7rftHjP8IzJAtZL1VuR1CckC0c0I7udh1bEzjButTnfrE+9d7PyF9l
E8N5zxL+84PNzUB1xBhLr1SV3FatqeP4fom/EiHiImws3kQbVHmKYTVy4+ytVCGWeuSvICX+tN5v
lbPohu6mqvBxdycKpPlnd3D3GkMcfpQo7KnUvlXa7z5Fnr1/5YKuOlGbSC2Gvs3sp96BLeOSi/Tv
k34UzR1zv/a5w2+u9PIlWE06PQfEiEIa4nWjm5vGHwKDfjfaUBTleq+S+uCBzjqC1QQbHSjFuCNd
KN7ZYpn9N4Q30aL7K4+uLfsWeqVmPqnXSqj92tZURTNfvY2p9g3PEabCKqBHiPOeie+WZKJJpLi5
82wgG2QZBsvpjRq3rZEMIQKy4jJnHH+v7PCW4DZ0x7b7DP6QlK1MSv7EQveI1eGOnw36830prL0l
DLfTODLVmjbK6oQSVRnpYNxCcOrfCN2vzPdVd1DlEXt4Vsdz4OJaPMZSgfevM0T9FDyGm9oY6Jgw
f0ekYnlbbA9bspEUbEgfURazhZo+Z5MvTrH4GxDrY04EVe9D475ptZBDMpWFFgLjdQIpLo8htv71
9g0cFhYrPx4Ha6tIO07bs3338oUz7WFypRxStB2NfTR9Oo5TX4V7QWHm0sd6dlq/bIRMdC8X4ehh
53UYw0z9iVdD3c+jPYttLCNUpW3RndL/GcR2rXwe3QwZVXYLRdLGwoRHQTJvQPvQlqXzBQWliFKA
GGZilUa44RYwexCS/CLJMgqi/V3pCy+FBtXNWqWzNJQxG5rVpZ+faEQIVEcihcsNUgS04axQ6u6/
oD2lum7MhN/7ERUgWUlWBpqiEYxKu1XBM9HL1+E7bp7dwsBWpRiGf+lnUuL3tst7hok+rG1+X+e0
pzOn1Uom79HMYPfsKt/XtamUnBy4xuFrsRPeFKWIqrF/8iec9EE4rGo8CGTgg/Pcj32yo+BM98Ha
+e5mz3TGWL8UhR8Wf+bTi5o/JWo6hsZFieB7VX80lG3mHDiwpOuSrdoGCArcy1VFQRg7w00/yb8h
ZEFT76LHQahRiql+2rPveA2jhs6qoEUJcpBmVV1l4vqQSCG80yjNGudNipIQM1A/c5r1CJrKNyFS
g5g2ZKGZyvA7thbVlFYy7DowKSMNd/LTP3uI+zuAnHBpMw3QZMXpcmct+tj54To0DYOOc0yFH9gM
Lxx3ibiUuaNOlVJ7HrxzD1fGLlyfpH8xTNQCDpOsCNJUWKkTkcO0iv5IeGH+jv4Frb7bcgRmAxty
Y0I+uSngY6tBNmUNZRza94TzoPI0DUMQXizexFzInWRxrhzDcAnFg2flPAR3zfWre7iXN6hhsb66
xmmgft7MLNRDSnIHfbctYfrG2d5jilwzMnMZNjDBpUaTQHrj2a9uhlzsEzqZksSAFdrUQYqQ73rn
4cArgJ9YbaoiIpzSipnZFhV+Rc9cUkhXd1DHXlq/noKqEWApNf0OpllND/GQ1lKGdjNTUs1RrQy+
n0QS22QPB38cS39BpHaWd0FLi1+56nJobj5WvN3BuoY++ke09Jg6b0iBaY5SOqkQAbswYUDX+9vS
DGAD1xExZ8WDrjCpLvrQVthLb3bv1TQYaIA3f59GraXa4TjaKRUQiAHDvtsS5omNIorIW4H3Y7Ac
/Sy9k+mwMGen6W551EqGFOaZouYw0iVZ6epPc+4xGHNfpkawlSFE06bKquLbw+XhhAMHrPRle6vf
TviBDS8CiWCp0QIF5TpfeYH4uUs67GJmUgkLrQBs0cIAGLyGaZDZCb6rUuYyHQgghGQ/9HL6H51e
7oCsx+7hjQ5Nec46LKLLRD0hJ/LbMouYTXDfielL2Mq9D/GZLCXrHgTKfw3hMUx+UTFpLIh/uJps
T/BOobmU9w86IxLaw5kYfK4ppIwkRxo0CkwYeGGAyxcGfMonn/NtVaZ5XQrDT2fdPw6iXvOIgaiV
FoKdCCJ8gZ6ZsSDeywdj5oyvpIneUq4eFgpoTrzG+Krv6n//xlG728+/YZlwcu7Vr5zYr+xR0rwZ
8Hsq6Ts4GyLF9RV0oAGlqqmV69aB7fdz5hpi+ZJK2N7oiMPVv4u4HQVF58wMq+f14gsFTU2xZVzY
sieNqE4B6TgbCIQZK4sa2ylHIA2CLnqB0QuLezZrlWL9j8ez0ep975QseS+c4fQ+XbPASiQp3AUk
x+deAcODebKeGSaqEYOkdAM+33ngW//oogBbutPT+L8t2qRVD5Y7TjA/GUno/1I+WAArj6IOroNx
NknEBueziH1JmwPb0yrkwpaE37/a8rCCeKW++jGx8N91x+XVuPLQRr8yqf0pZqkqhJEHmgalN317
uNGEeljC8sKGAu0vWdKfTVX7+YoOItBa9VnCQW7+oUBBYD9VyTdGEo9Vyl9oNLeuuZuMosYBnjGb
6P9TpRhIvWjw1md0m+twsdWOY7jTrHtKa3l5elEhMreHTk6GBmEU/zGtnbxJ9fazrLuHLlm9LciK
w639TrFy9l91ln7N59zjvWGXhRjOEqvEcMWO5GcUjrbKak1P9K+RoF6iU025xBYvkNTbUdGlGBMU
mhH4PMhDkx0YUTQGDFnDATp/TBY/hzDLSkwCYlJO0tvxiCK/PAGlmSlBvvgivKEyHOu0fCMViAi5
v6puVrdaRa7NokuNo+AIYKg/RDQ12aSHxRWzbhXGhcEpk/PEGZKpZUL9vhlgmIUVpff4kmWfBdku
7Pi9cCr5gUPbeHMZMl7U3T44XRf+aiO9hAoeJE3RiQm/jWDVyJKx6SMM6Coacxx3vNM2ARhR17Y1
tZfgdqxLTjWfyGf3GKZi4HzGqFDvUhpXm1dkyOq9ixyxVrLFh0vfsmWz0Z6qcHCxf5sVEfi/oUss
1DW336vXk8LDv3CZZ6E60cxStIIscKKni/0OB2ejdLoiXhMPbOWFDsD6T8bORXkuEu4bru7cgLo+
AgwOrFF373Cmzb5gm1NKHpbF0XP+lkqrUTJfxNIY20zUkNALtb66248sRESgGQL//3bXcYUVZBR8
7CrDEiVmx0F60OWnnyioPug0UWwLYLr6zFZMy6hfTKg58UxHfaQLpYSgm0tW9xP34z8AleuDLQxg
z7NAvzU9VuKLUEzaEQR7mmsN/IrsxRbgxPFpXodSRdHxi7G1BOMTSpLotrIr70grQsRR8mkLw0v1
62qNwt35f9wsW3NfAkiHbMUozwumYszMq291VdiQdvB/EQ7Z7igLkJZfTxNL3abkWYiqF7LnKx1T
dSlTbleuA7Brlnj690QCAju8cZW/D6eJK9Q++4wT0NMI0aNsm60RfpzocJj2HBoYoAHhSb4TD9tq
rk6L/GjqwGXZNBBANVVdni+qIucNq3b8tCwhSEnW20j97v9SyuRNPG6kJH5ZvZW8zH47ZzxgK7eP
Dd++nrW/bdyayKPeldBF/4E32+UG/TOeh0h2VeDjl6VnLjjd5G6OdQtKwN9QBt1+8BWxgevSQ45Z
DXQ+LnoOKFdJwtwJbz6VOqrKc0S1y9XUbJ9ggDkOsC97YD6VyCQh9ByF6PTDZeonnGUNIPrHuVkS
OexAb8/0A0hqv8TfMkOswZgFfLWNPT/11L+1z45VFZpPPr2vO9FqDz1FfV9utU0h9ib5vaYRc1Wi
Z1JxAFwHjxxdr+/6nSXDR5vTo7CQNMxXbqyznykDRZG8gyySXdHisAHYABI+Mi7GKBxddLUdwvTK
sYeQgZzOm+vFv/IbDBg4/TAqqQro0qcwi/HQQE3he6/tgjvHU5LNit0QYob8POByO1s3Dj3uHrXm
zzfISYcNcaOFnC6q//T03apy1AGzzdmJJjd7m5Djf9OwcBO6c/zDzAhn21bYhzRtdhbvVQOv1sY7
V3WlP4JiZx1pfWlo9avyO3aLgnJp1I6qESmGsCYOH3MAA2xC7kR9ZZj21Ci6kB4TcahKLlpJN9zD
TATZ2nKnw7y19WzqUoSE7Xj0Bc2EDw9IyW2ups9/Oe0/XJ8c/8fTrrhJ8WxhNGFuH9bYRZmUARqA
iANk2QMPaC3JsudaXJvb+gRJr/ViVq1hOvJsIOdBL3kIuBDqBgPiHi9jEdWBX+SsgN9GGNU2ZBku
HRZcKoO0TcVhj9kZhVRZsqMqEKkh0SheufDypbZM9CbkxKBSY05X+YIXWfRWTsI62Md+NkbjHDK/
81EeIZnNpmXlH9a4E/690d+VNdGaz+aMHtENiKCobx2xr2x7S8LiKRpEu0mOR/NRaAmpb++ghpeY
MTu40PcQqoyDhNbYSpDd+bVIDbP2uDgetyILscEa1Ah3h3lwHGQai9oyFykB/2NiOUdxEPCO+sM5
Qtb3S4L52p+wa/n2odHBlt0o+jKSHgZpxkaMzle0ByuzwA1s+Hu6uiQxBxJgnKO6t9GBHM+m8nnv
xqg92mPSCJ7/NaFkU3/USSq1/7cTgh534Memj/iLHFGoB9hIvaEmsnb92OAdj+NZPQbyfUxrmS4X
AmeXoKqvppPKeSNic/gew/vWx6457d1mq9zLnFhxngJNqNAqK09UP8ehUOz68FkpNrczI7AAkDvc
U6uNWzYNUO6+nqh/MRkf2pJJZcrmAPwK6hfbXK+xLUwkM+0Jl7FyDUTZDGFbHn0fRnSrH9sIys/u
3LAGvMYJRR016V43K0NoLnSKhG/c4KaZhz9EXeBTxfJX/ypGUm3Ulql5TsIJ1MkSrZUBkEIuyZtB
XefVEQC/vz24IuJZYWscpX57ko/35wvZcmMnfL7IYDs+xpbZoFuF+nOOkjYrXC2/D7dsyM1wH3Q9
/Ze0VQthbNtL5qIsqfY8fMoFqJokDQt45hgvMO4cakcp27hlkUYeOq/IPXyjewXiBxlbSh/hjtHh
PLgCldQOIVlPk5AruONCBcZc+TaF5dPLU05Dk1g2HWUkbr7b+ct2emrO/QmvlZGGJRL71SR6t2Zd
7UuuU9utQENdOrDBo34RITrG1ff5ndLQOxNEAbxA7f9GJXksRFIaQcnMGETACsF8HAmpPpH4LB0A
LevYDeF9wSrNDCBJl+84tXsfDVsXMDmh7clmeVXjLebU0mHss6IxkVsy/RrvbBTupaQ1Qeio5UJT
t0bgG6abcrlHWMpeSai0Di6+Wy7HS1p2+UmX+fv3r0ZwF9LEHOtMsVgIvnJzsO905q1feUtG3apf
XRaPK3zbJXZZVBMbTvEKmRDhTM8YGMxZUGzmaAZauFCD+3oNIWR+99QrJzsAmFo7M6NZc7t1zffQ
60SqW0offN78z0lNV7p9U76dLKDElRUtYGt0QzTokPHqWXrC23gLz8dvmnSgTsNvM6fVgsPIwXEe
e6SLJ/k+hN3YOtyuM5fsLexf/ueQmygb/OBnkXTjAgXJhTnhEZSNTZ7+IfIGs8Bu1VhLaoR44Xfb
NX/pKj3SWiHTshyXVp3ZnO7S73qP7q2ip8I9DECFaHmtwO+9K063gC9NW5IGJrG2kmUO2bjvRAUq
pe4A+FWTBYDy3GuWGRQ1VGpj8VBM1jjhEh7dfg7zA2rUk72jjcHWK/gZj06JnmGBwT/HA45U6B89
UfivwKogZNVi4s2Eoab8WFKjswS/ojkXBWx4hdOXjyo4bVqW7i4lR/ADIzeCp9pdsWas1CyP/3p/
i76jS3Cz0yiHJ/rFcYu1cDdLLQO9mF8phd59UbB5yfkCgRgD5VECnKvQJ/3iDpyuEkdAdofQOjMX
g6iCHUlTeuYDurwCNaOsUNqXS1lILq7lUCdOVgckqTMOgcWaxRdo+X4elK8euAFgsJv2wKDyv3tJ
bbRlfyucftvEP+PSjbO+GAfMQWT1peLcKKpi7+OgZTg5/73BwwQJ/hy7WfYgy8YGavZulgYDZSwt
fOHRqazaLlPvzl17UseX6OJylgLiwinGokr4jQSlEL7rW/8vS86zIn2qSJC9gyP6aXEk6ZMQ4+KF
iMdTixt8q84hfC1p3AQviJRhgvpgRyt5a4n7bvW4yUPSVzm6sNZiPiKIl1Xz5fNLesFJXwMJh4eo
M6UMW97xpJyaA8ScD035LSJoMoYRLhQo3EtwdXfmtKFjo8RoS+6YZkYLbo5MfnbmMmFDIJeQ8cH8
FrpF1FMNP6enfw5bArVB43OzpTGjaKnFC73LMGVLWBnOX2hipys2UYo29+MkwKxES5o8z0/AXDAh
hHUbKwCgwVRQy8Ckui227sT4w7EF1/ij4EY9nCdLmGgFnd7/eOyRTKCKIICbcRgAWDRNZfcxBkYH
3SCDiDoXfJYy+6lOovWleemwYpcvLDLOM7jWaQexBbVcyYJpASqKOA1vENokmFcG2UW/K/toRkQy
YmyPHPBjphxiBKgMx5c4BQmwmby9nMiQMgbPhRkZJSQC3mHv/GawwstcOD2KJ88tzJMslr3rYJR9
k3ihuEzoG5trN0Zu3ADQlk6vw+n4YET0mg30Kwhh7cShbl+4uNClF+dZKboe6Tosqs3IOwsjhCpB
ZK+uQXuuou6SvrSHXH3RTcB2W+TJONu5mJN4UzrfQgHnzkfo7V3PV3LQ0JSYOjgCs5rav3Zw7gcR
NO6VAAbA3Vlm391nIgXo2TFhn+89x9KgwD/yp3XKZDMEc61nc3Le8czcoldUw7x+Iigw4fVx9b71
PaVgR9TUKWUNI19Va6qtQgPnJrXGs18EAAPHWEaPa+iVBEmkwQs+CCmMn1F1b6WmFnENOJJy0+ZV
QyBp+lWHMyuGWzYfa/NFGGHpm1ChNat4XFnqZ0IJaViFGcDJxsCiVurpRBPkT2GyBQiC2SC28YKF
Vus3/qw43t4Ky63Q9o6lD2GnX7aJDB4JMLKzmocVvdstRcY1D2kOhD0v08oXd8XEkOVmnYLLGuo9
ikyjZ8qBbmNq+qm6x5g3X6Koa2SneKGiQepQRURLJpWhUkzpnCnYIZwRBAAMaHgT0j3O4nUMCoDX
KuFWskaIIor9f0kCoQ0OY8cVYjDrk51Ql6pg8K7Z7GNC2xgNixYI39iKsImoKbpQUWoivg+lO3QN
aRqhfOxV7b4CmajPE+ioFig9ddDn9caGeMwDBfbrTUlBxooatw4M8C/lzQ4WvbXRmpzLvYSqBbxs
wL+zlJRrs7VYarsN8orYuPfqD4mCLCft2afNbbrJV0WaYf6LM5T+ZgmZ/t50P5jm81144GId+j2z
h+jUcaB+FGooAKhQD3UfP3AQ2JzQPRLcy/UgGI1H8H0N7/Uu2XDUYWjDj0+q5VXgJAJar7XOPBuV
9Bd4Ib0I+LnR4xJPQ/HKdD02x1/XqLs5/lPE+cLxH+p2lD782yFm08lAq5XQuYtCcY5gFZWeTSoS
EzdRBRzrm1unw04ZVXyDRz6eeN9fiQQbexYv3MQerFtgfMkknuMHjKfcxNsnq7OQd1XFM11glNnb
kus511s5GGuocJqvz/jZx955wbgfGO071c6kT8xxWyaGyrbLdAdaB26wWFVZAG9b3ZwkpaCJXvK8
kvYujNOPUojTCjn7x8I2VxxNQdZtrhtgHv0+PdBSjergIKrkJjiA8E94f96Z0wQFkjBNu263cAHM
kbyIDjnBYx74JvhJXb05jem2NwdLOIkR3JeuU+XEb51TS79x8R4UE28uw8KNsfPrlNb0om6l2XVQ
Ekib/49cWJjV5xXyfFv6Kiygh9Yd/Nqbf604bJcxQ7e3chrdMOn9N6zklhsmGNkVRUwcX60fDNeW
IdJf1O51zSmLLRbt3l2xIhgWJu9qLIS4ZcxuVu9q5vF7QG/zrBu/UooF6EI+KUE0bkQ1khgkvHPD
GYZI4hoUSab6p3z2nasIJ1vjx6PTnlteVLU/61mkx61Fr4yWOc2Z9EEyFV8AY5hDQG3Neq7ko3wS
maNjoTup/2nuuMSxVM5SF+bJi07uy2FuGlEmGt/wWhNyODHu2MjBEW29BDVZ6qQurk7vmSokl+uH
PYoorRI0KOi2UViRLTltrgwrPy+/ZT0sgrlQ0DJ4QY6mmJw+iDKep/1pZz60On7/V4ZiACC/m/lB
PBU5ZTHzdUqXcaSRy98kEqGzKAmIB3vdUuyGoxqiJV+okt0fXCwWwZ08eLNxNLY/VtrzFCgOy2SU
YD0Q/69fmKg4lvOZQc+mYOsBplngPihSHm26WY2OnCHFx0pLjJoT0TRoKt4Dv0HMZh+HdKsuNE5o
nO4IZZnGj5OibRF/c8BeI9thgaUy6D+foNziYtS6Dw8x8q5asnRyzIhccc/v1SZ6ebS3eFEf16fw
awPXIfzPK5VpmDy6R+DzBqfRUtEyw77zjSqJB7pRtFUfb7fRqFqofe6KoG3cExEDDYQAioyp5T2M
7KZsBf3TMT8aGeha4MBQTojZeqnW3AZ5wnRFFt38plgEBapOMdZ+mvIH3nfUQUncilk0a7Pyeg/X
FM/8ZeaudMWdhTowi5EcLvQXU04mXPbGzfo1ZRnpARbpn23bApcAXGL7gQmBrzj82MDXrC6IybA8
zB7SWCDWWj69XixpAeN5WmJY8A2NyULHL+EvOgsFSn7uNFJhVT/t59BoAEhaXGr185+DZebR5k5u
Zfcpsg/NukXj4SsZ8NJr5MmJokQrpyIQJdNciyGCcTx61gQ+OiKDIwqKt+UFA48zStG8F8QS5wqz
3ZsFXgCHCvGHhDPZRxEDiRnf/4/PxD/bYA+V5iuSMWYNCjJ3iL0LgzlnUNwIen180cz21U0UDLP9
e81TfEYjxFRq0ulP8F4RE1sQ/3xKl3Us+HO1XGyVKQrcjafDUDJvK770BylihkNGZp7TzBHQncQ1
9PynY5RW07pnA7sFwdUwFNQ1A2Jq3Eh/2xuSKq51BMLGtqvUzqc6izguzVOAQzFewal3gaLciZBC
NFzZNxqWMc8GpB5a1jo1bxHcRXribpvjTUIhFr74j1hEkPAvh9aLuK2Fo2JpWwmElkmr6ea4c3tO
1B3uKQc3LBgdBe9wha+MNcDCHlgEX4byB75+AVByvlrPU6eRw8oBxbKOVPZRBpLf2WzYJzsPdTBt
NZrgYc67eUne5/5EvMyxunvU2F3M4QeneWZTPgI+XfZOZgv44wRVHQyfcv8qzYrykcA46Z5wVVYr
nl+q6iP/JNPFUxZawRytqhIGG+8io81XGthd7DF9xjkZSkGvzA8VF8YlE62aoJL1Tric5GuFCx+j
X66KUCXIUhs/+gbiQ2xaA1sT1D/t9IVWZfPbPONLGL4G1ruOz058ed5DGqxPAP4RTO8Xd9MJ5M2n
n56lIl9ztp+ldeI4K6bFvpOnv4Ttw4d5bL8hKWoqDROEvc6IEOD0afZIGRdTnqf1xP8fRORqtsA8
wmdgKuksd5TaqB04ZK99IwBt6RkQugln5Y9rzhv1p20Rvbl0tDe1oVaO8GYWbhIltwAENxmOXdpn
lqPeAU1hAOupk6hRfrUBsUxtYZsua4CTdc8/xrLi24bl2uoTsP8EfbA9iPuiSBmdjQzBPEav4Eoc
Bag0Tsi39wwlHXg99hb60/xFHCM8k7/hpRcywkPvTSDU1rtObMX8Sitlp/JlG4EP50eyTzVj+F2+
36wuyKP4MiL+nvj+jvhyqP5EuRa5OTodIMpvZk8FAqy2+3URa81k5MyLL2qdreoF3ysyUVraE07z
My6t9F1LDxihqWv7EDst1Kqfe/f/ioqMK1S7ECkV7KRvgnDIMmT91yGVLcVD6/2kEDp0DHvw04La
o5WJX1qPTMNy89JiQa+J9VUJqi3WriIeQR1FuABOMhMFSpKZZP23m7a87NBcPuJQPgFIF9NZ7BUF
atfF+y/Rr6zAYYsb1LQMjQxQsRPNTutLOE84eiUJ1kzeqaGDdW3mq0BvPcCz/U75Otw0fpRn/bxp
AO+hqdlbF8wH5ndXZ5NZi30BbM7PP+X2y8tTUtS2nbPUJC4bYgsC22d8gM16fVCVkFF88eooN03V
ZiHgmCgEM9q/GwTDrFYjU0XQhEo0LFxVXmT5/IXCWerlYv02b8+MACFtIqKX+9uFvOQEYQWw1VyJ
Tc642s/FuOFvtkAyMRNtnG4RImKBg21FjDOXwMbEptLvammw7LoyFU3zJM5bZINJkwG5KUdezWj6
w4wZqbt18J0lpjhN3yqj08iUAYwsKzF7QcuDgCv+PSVQEZWWToyh/HVMP+zjK+hm1COEXWf3Tuj/
SQ/umyAQNI/UsTK/f7k3znhD0/Kdjd2O95/P5d3zqkSp/YuYWrRRtqqHWPzWwZTntGpuixsGidop
32DqczN4x5PFP7zZevkvnypxtwJ//Uyg07jIkeSuF9QP5UlXcYBpg5as+gcda+JzErPZAuf/ll6n
fKOOg6B6TS/UPCLteJHQzDql3n1eLHZ3ng/rBEtrJaYia3ZfbHvAOXroIGFOA5kKpKWiu/W1V4uS
/vw60ZYH8fI/alOhHDQSdxuMaqVwZijmuJc/5IZ5FEXMCjQz6z9A6ooMAJMJMUUVzsyKxvI1AX8M
6ncdnjhZatnQ0cXvFGCO+gRRccNpjG2q+bMl9tGaS3tG55LVuMvPCJAKpApufdfFLZ4UiTfEGjsH
i0wxf0nYs+BiRUIFzQN3lDQdpkm6F5LmeTzQn+IA3nCIVIH3V999m6DTU9GIDgv+LbtycyGFlg22
0Jg9CMW24m9gCfUJrk2NzrfXDG/Vg2N+h1VEH/ZYmedJOSnkHXrOZmZRd7fWb5B/PPoqNlwBb8la
PWhH/n5ZN5gEDlDwT1N4aMgUiuRP4iBu5ywEf1zfUITt6pzWkkAseQg3UERtbf1DeJIBvYITFxD7
ghenXT2knMSv9kHNBb9RWKZg01rDKFqr8xlvdfL4sP95CTvLKwodJtfaywx0o8A6LuvWRllOjGAW
W7H5KfpaqJ8bYaD+drFnuObCf+EM/sCJutvtJkvp0LcFlXU2aD1r20GhF9SGmkRU0kht4jQ9VaZi
qzBeS9Oi3Q9fnihOVHojtjDtd/ZNIef9inscM68I5sGRu1JjM62fgvkZ8s2JPY/qbLAVwvEIeL9O
+edAqzcat4XBDLjurmbaVpIDqjfnOIBqXOA5osq9hqq50+Gklu7u/qn3JDUaz2f2aU/pDRTWXV33
/k+S4qLTqpfbgEbuaNY8K37WqScLuTgAsWsC6zz3P6maAF9Pyra5/oHGtxR9lkznzvzyxcrDMU55
9sTlT/H2ZAb97rjyNVO8eXw0zsL9oAkVpFn7osQ2Y8iNR1vBrf/CRqxE9PnUQf5+bcaU2rga0ytB
o7iRj8JyXK7JyVoSq35Hxf/hu0MSFcyETJ13/Nrjf09wwxAwDwraojIVsFKoovzUTJxDDoCy94BD
HKOZT8l+eNxf/flvO4FWU7ZPMincY/me9WR9qJzek3i5f9/65QBBo1+UMo3TE9avqhPAicNrR6rS
yMsnheXpJHdk1taMx/5DPNSkTYE+grUzHyT24vGuravsdw0lHgqvBFxIizONUmoYiI7Zo2b4OQqx
fvjFRplr97ORXG95yQBVHuQZJ8WNP2+WyyyPIE9DNoW3jh91QiHQ8TngIydc7eZZQgmGdgrel+xR
hxYN/iWcWl+WaqAyneAp5b8oCf7wdt8CrYA9Kkdf6sqOTCw1qKh5YvYAwY7EbPdukswnnGTvjdzA
v/+ZaZMOO40u41bznG4p/+vM8oVUEJD2abGoQ/VFQk4XhAI9O/a+29Vsr2hyQ3Gw69myzH2GKM1G
+ogUkIbY4yUvijiLzE05nE3idgMJ/IVZDKmkvFKXCfjGlPx73sG0EB+MXqpWpOww1nhge3/sWi6Z
rZUuiTlksTKlYmu7E85kRugnPEoQWTGgWJq9s4hAxyV1JRz0eBaBH6uOnwbXphY4UXc5rQUkIiHh
CDrJev53qV6Sku0ywYiUNrSn7RcrWTCEJWobI8Z4kN1+62PmcUvhSAPk36GFbv+De0jJDZBnHnnx
PeIJui0Rg8AMdLHGJmyd3/LlFE4cW06ab2081vbV2ZMPdmmiVhlspbOGAwEE33/pVDJqYdTZHZ9R
MxfOannVPoOqTXdrynMduDWQf8Z202O4A86foXqwhMD1ukvpz2UBnskG9R1x8wpDGxMEYvBPHQrQ
fDzD3rGQoZhXftvr4Ayuz8E42NWIUil/2nb2KffVdJlFjIlgXUYjCd/FumXQnty1Az/x6Msr1GFW
SittwSbAfMhV1j3g+TPMfwDfKndm6RF4pcuZ53/tRAis3u36OamHlSwJFxgo7dSjuRMmLdlcnCRO
SYdkkCheR/MshYzOIrXNPdyvbTR4JSx/aqEJZlWp6sECBQfHdqhk8CJCwDp0iXA+XkGovu+LiG+D
vS3ALlRwgSEzqWAQK5h1G+ODTNcZQosMoN8ce1bzPMOEDYAbouh/o3/JEH1zt12alGb24cXuA7ht
59krdCQr5MDRONLH6Idj3v8pz95UfdwZDNzo4xrbZrvqVTYdEiBO+bIweLqzgKAwiucG7+/gmi7N
1fxkDKmOJuK+nL4t0rpIvq3RFLAhjzOxVGi6ewBGher13+WEZr740EAFk9isJodZmKBNrVqQsrUd
k8pc1L/SPqSpYGlRfsuaKkElxA2QnLQ/9/TExJzhC8cAN1Qq5xme+2XnaoDFZ0eQmZeukG1m402U
f697Kh8rKfRAWVvwOkvfwxZg2BP00lfUvb6KBmoRysKlHXgopUIpf4oj8u5T4riO/H63f9ibjVTV
Hts97AYF4E8Hyja+a5YEODNdV+1lvjgj5wZvtPKooIRkDjXXTd+5TyBNgNDswrjqUKRhZr1Xy9Jc
Ykso2AVdIULUrNI2Lz/XVkP8Q1RZgvxTX1tNRYDtWJVwMJ9+h7urGYFLWt0HmQMFEVZcTSb++5kj
WZZihlRbExewdTBuKsfqit4qDK3Apw/cSF0ZQpB+z6KYQipCJ8wEyvnH80eTo0gVIAOsLQY+uOcA
S1L5YXrh1j0iPYj+1yWyAeeHfuPWk7G1Bvw7unLCnNwEuLBTBAQl3Jjrnx/IGLuDOjqWmI/Pk1FW
iXwi1u/bhUizbZWmpXMjeLNdglX7Z2pNHuDIZmQhoFIFzu5I046iAZjmpwsR0gcy0Uj2gZONaBSE
JfUKYClXYJGaYp8WwuPJMHmic9HYlwamquos3CjMHK9yelix0T3eYwDfppondLVRvhkk7Zk1fWlu
g0LKEkGTWECuefZMWljYvj7E+ME/o6QIhNO/6zCgrqJjlIsX+ovbpS/6zXkCQYjigelaQtwHv16n
NAYKgRlR2bjd/nCqXGrGpBfNKODR/im48Myw8a2AfxU/T49fvLF5siTFlsoc3F91MLUaPv1600S6
Jw/wneDcLRJv7q6bvGKWA4i1JeqHpqtc/SyfK5uG34ta2JK3QF97HqgEtIUhy3L/MGlaE6h+wcIJ
EWHXpmqHM9qBFbSRlJ5nJp9p/OlqkQGcqQEw50F7TOO6TUlq7CerJBh2vs2CO55OrHu0t5Yw+nAI
mpzPRLqD1Rve7qveR1seLq6jGQI6KVYtn/hGr7jvXU3Q1S89Moe0zzkP86625RWoSeh60ZUq5z9C
sx7xwaTTSPiAITD9IM1xpulF9yOlSymQICJ8EOVik5ThzTHB5ei/0qX1fpbeRH2+4RX5PEv870XR
ZerRoAgIV8lvZ9Auow80Ga18jawTOqc5/ktv+GVTju03YZd+D+FJe6nQK4FqwwbLN+O2r5IPObxn
8SpbJUDASoK2zbtKjw0TVptoHrOHMtvMuMSBKLuT5jUGJAeoeoDSoKAmNXsDmd4n9Zgtes5+99of
3hesj7Lq12nGcW0fKsg4NaO1QNlkwC9Y/1tFKxMw7YX6aM+BQGJBJa7Y+/26i/p0nwVj/mmc0gnz
PiBOKh5tZtPEHc+B0kkN+XasdiEdZrr8JBXJamtavk7RDdHD5/tNOewcNPkRrZYSdmbwVNR/MpRG
gdOu+Kl+wxCItYQnQTcH4w6j4pmUjR+aiObC/mlI3nLXn8xxpeCkT+tpHGE8LZqetIRh7z4FdFUq
tdAl523Yv8mJHTIb/1fLMKQqnUTCFeEy2r6FRfWYqW1KWppVs6sEgtmxiDJIa+ma9RLfUeoLZ3OZ
hBu0KdQ0fyk/ZKNKMH4wCAtgCIqsoivCQXG0JCbUNJEs0pheAuayCDZwHtVwRyBY7w+zbkdFpEQv
zptX6yMNS/7ZC+HjcV8j3GNrolcbYJHb748kn7bqBq0/mwNld4dLEnpWRACjv5n8yTZWUKHt5B3X
u93Jud8fyvnmWlDvXK9wxTQKVQoWsSd3zmjMiHBdsdMwB5ql530WmxoNTN+qGocCgoSpdgcGqj+K
NBkJdiZoHM9bDdv2AA3jZ4CS6r9Lsqge10wZhKWRtJDRHfiA0BzOTJMXfGRET2cAoRF+OS4JWMkV
idR20ufal5HHnZ7N838sDnFibgNauw/GSOZaZu0/2FDuXNG1mnoevMRXKAP2RwM2ePf+y0PGip7V
nrY0k4UBjvQRIGpbXYKm8NF80JC3f7IDS/Tafs+4cg68BRRLr8OgW0a7D3rxPczMr5W5KsM/ezWT
FRfVYFrEKEx8x4am4yHcbfL1t3K53LcLwOWrE2ZruZYIHJCUCuuV38Fzb3nlf33d4A6VwpZhYsjG
QLdisz4sno6yKHzr+7FZDBaI+odKXs1lMfEwHeHnOaSXAL7fz4e9xc+ffwdgsUc+wePrHeXq+rQg
Qbi3xbcsc1VTjrGwtjRHHxPl/mbWjevJJfTxk+lIIFB0cvT7X5FYySNVqhM/H4D0L3j8PjQhse1y
RTlxKBOAWVwMrp0LVDYKNcXqtyIzz3yg5WN5OcJMSSI80JSkaLnuTNMmC9gg4SvtLMZkxt6tdqXZ
tbg2+80n6xdw7MRYr1uPjhRNt7PiclxwJrKB18HUGq/Jok6uYxmDvTa6aQhMO2jBCEVqBB9H2MQm
TnDc6iM351DBM6CuqMpQyaTn1ln7xjIUQ90Ho35uC50BxzidYfa31GuU/Ln5MMKP30h0+vJMBvvf
BDWGOD8d+/5Z5wvOFAj+bblBmNlvBWBtN0VctNkQh/2RbSMH1DPHmbJY/4Cy/iJOjEUxUyIY+H9t
xvVdAQGCjgo2/Och3mF0VPn/mOr7xoXW7LvLZYCvJ6/mdf8bQVvRbzvcxtUIfPaHlxp9nm4nbZTL
h5hM7uAF95QJWMr+L1yKshlFjRi+kw/TXRS/krpxquyq87btxWbyBgoCaxDFita10PdOt+m/X+4u
iDo/RW3enYHu6+e2r4JUr0qcfEAW+FA3UcIJUJai9P3ylmyBcdooiGtcmacWsg1WMAwT5eukG1Wp
30nDcGBH6NAvSNxVhULs/Ksz+8GuVNwhZbfPztLVyl52LQQ8oeVl8OpzSJZZ6v7AdIiw645WReAw
TSXKnN2UPF1s+DUIBg8eykvD3aQ6p26YEp7XziLmFWwT0Fiz4hJ4dqdZwClLTrEp1pOilcUgmJbd
SxeyvPPT2cthUAxAA+7bHQEwL4c77BMuJHHU3ezZE8r5nUhbJNKNUgc8eGG7z5EvdtXJtSO560AE
+h4KKinAZanEyPBfDQ6uJ71zX87hGnjiEQ9rQXhbxfN0MHrW7rDtY3beKSs/W+sM6MPDm4axOmul
AH2rJfEB8ZOcxUoBh9Fw5Mv3MsrlpxoxsKX0NoSJ61Tf6kwS6A4iI3FJUYB7mVOFbytO3SRSnX8Q
KwXC2mtZNdSb2Sf2oYuiZNLxol/qaNx9hSk1e0itX7f+3M1rCKrHKMGoAfvD3svOIyF1YBRZlKlM
xGWyBh/KUuyCNgWXWF5A9ew5H6etdlJfnYCEU5MZFkEPU2/jzVarNUHQx7IFRaJZISWVNqJ+aIvH
pKL2CHA9gxGPwrwZxS3SqAC9MduEEXhEeW94dMewzdXuf1D8Rx3XjZ8dgQzvSLSca5Kb+9dMFND+
ggTYwFjwCFm/wxw2y+c1rrVtPA3Qf6vTZAKww3Qb1dVZPganeqTOweODrQse2xAfRSBOebWYfwkZ
cnHAfhRc2sHMOmFGZgXK364vKBRych7K5MtbhPqioULdAqmdBpE/5FFTRDOVNypUeg/tsEom5AZc
Rk15XDhYPvwZCBpB9tCtDJAL5FFKYzyCc9ywgLC86ykNHqLYZyRQJoika7l47BQJBaeZQayE/3fL
jUQNARkbPrVPXnWKS+Ofg04Q2DXeOC0z7NhwhJQn0jovdXB5rmEOJcgZR2qymTrVgBkAOIDr+wnq
6+YMsUuw1iGEa77Ht5eC5sniQ4wEs/IMaFsqtboBnb0eO+846Gq8t6aW5vIi/SqiM5SNafHCldqC
//Rfn/rZY/XQgzwxRVZv2d+Mm/+TTwkzCx7rcOBfcnx1DF/FMQN7aGZoeqaRy0VRB0LNzrzPohUm
OZ4IaRl0mDm4IxrtGwUStD73WzKo397X1Uy2AXefoWSE2so9oPfCbc5zWrTI0lZt9TWofyvOeIhm
QoEbD0BYeV2eItusu/X7p0sEUuTHjB5SqXHt6TwI88za7Qnh+NSAfNNuxwhMw1fAsCeYeNctU09y
dvmIkCtgWdZGNZKY+UA66dttjqidiw6J/8ZadyaNWU7waeETG7rzW7bEbqmYFwCxJDYZIaS55jCi
BalxiHXWT7o73QUHunmO11ThRk25Exy33PnKpG/sKTemAHyzIzDP2jeV8VYTzzDPoy9RK2NBAYQu
4/DcIi1msvGrSZ5F+z8S6dmUSeSsT/tJ80msxrZQGGPCfzBWuOWBuIaEloHMMl/6jGPfiv7cVms8
zB2Ze0Rlr2SqU/0+sKaD79jhoFnUhyajZepnWN+LhSIrVZneodQH4mCrKibHuK1gwecS7O2qVg9X
E8zE4XOwYGVWc67i2Lh9YEdmVTqeJ0WqsBq2yzHr4umlsJ8rglRSellwLeOE9zaf5b9WUtfFVkNp
sD8gDupNzANnfLMes9+pnK0FIowgtLShsr/zklEi1voTvJGCFc23wO0+doja4WD+DkGCu92MaRFw
Vnjv/VmgtSthrNP8wci0Y4cX4BZV5KzkJEtQK9uHy3A8tJOgxdgNZACXgECtnv6bafRjqNYf+Ixx
itgmV8s0BrjasVolCunP8Nj/V9dAiZ2P0kWrJWE/W+w+c4Otu8iBhKFUdD9WMpPRdTnb5YfhXTUd
icmN2SoMPNuYsSEsO8TxzB1Sde8oBLrRyS1OVfybIjRS3axvINGo9TCc4tz0df9XKNAEaFjmyY/d
/6yZPLOEo2cgb2lPbYyoqdEzmFXprdzmGGRvHhIgB3zuGuiA1tBFvqDP9C3s242bfKIwroTYYR5n
sCbJ0DTedERwbc8FvDzdz6y4iRRHDwbImASKd5u5W/KrvebLYWDHzTQAdoF80SOONRD+p9/rxzqE
n75QCUL8jPPgGjDh/Ze8ro4TY2wQqEnXkGrlG/LKMILnSqM70QpAl+MSIYEdnbv7xC8BfHHCfIdM
LbF7ekBzZTTtsb1UhQyJ32DLtShtlqLZauNfhM2B7/I69a/QR7Hjl9MHAdnfActc6SxfCXAorFj0
YqytCmzvc8l/I33wDgKItOKNG5GUdUV9yTS3PmM3YRjlg5Qh/wqIac8cBNXmXQzwtfblXUXzca5N
eaLJVtSwwidVqb+J+y2OaMPvA/4GCXdyZjejDLhbrD3/3hl8TJTDNO2O2IrCwfCjGjP1lbCxKMVe
WWTID+GAtzUTyFJbHIBV05i+p0w92iDM/g/YmnkL4iGgrTkUqDtOkxGzydh136FvsnRTk7uAE3F2
dOkyvzL8l9gKpUB5oPoKfQX29b6d9RMmDbB216oRkjjCuJ8AQKfS92GxUaZ44/pO3Zb5aMNSfrgW
/bphDoTv2F7EEEqBs1m7/dZGo7cRnYkrAOe0qQZU26NqX3XzAusAcSzcda1ZMQ1DMyIb1K/eLTTD
75lkNeXek9Is6rshhwXQWZjnFZhA2lihGbPDrx7YN1ncA/ZEOFIOx29MQGTWV4DdjUJfCnYBQlSe
At/gInT+mUwy4uLUrQA5uejmXpRIL6QEAJVfNH+MxpPZB4ceO2k+rcz0qJ8IwUE7hccHzrtHG20v
I5HXG86OqrDdhAbJ43MF07bW+pcQQLiKSPpYYBZX+TGP0ZZCxm4gC72+96JAInOAMry5Z8vHEuvS
sjaaZ1fb0IP3wJbMN1yXXpru0hI1QXU87gIKoSCfqrobE5fE2gBS6i6phUmAYD2zyyL6rqpuyFW2
EpKm6YDIXgVwDhXFPDdk2ePTMs1wOPdRZ/tgkmbn/JgkzT75Q7ocqMe7qYC2uaFfeuBPdDV0bOgw
eKzAefR8g4l6q2JWuAY8E9ve6YhizQAM0EmHwMC38CAN/c3/en/NZHqXwcXVzaOa79cvuGwXXF5d
QdmLExfS4eVh785cXmiTO9M/6fswxxlwgkptNO14FavOZgYtWOcvRPwe+2XAm0oFXn21xBiouqim
Oi+uB/IEYItTxVPDGmC4XAUZ44m8/XHLmberfWdKcOEpaVEye+Ev7N6/tc9utIXaMsD6tpdzVNOf
SH7ZBuRvvlxfSP2fzugLc0IDLjGjl0cla/O8Zq/YfamTc/KU2gv5VIP0cvKUlw25xC9Sk3V0gvCr
+Kbh6M6Q8dVWTIMEPs66goRbv1cJOe9W9nF9JKlgu2AmpKZXQ5exV7EHFXnPvwJfhOG58OYQeg3l
0WvDxf8TWf0zP0+VAbLawp2EL5mR2Ok6ZL3fYTrO+nxiG7E+Ep2tGT4QgedC43qoqj/sFXzr0r3Z
S4fULbvee7cCOFtcKfIFSkZRkZBp4F5Dk/FDYM5BBTaAvLBJWd8CGOLcKTAO2GrLK6PRJkEYnIc6
CWzwo9GfR2rzfOYwKf5va31edyhGZYy9tpRyENmrdqPEiNJGKwe3Dh6R6uzChGLMcjAW23IDOdZ2
iMmDY4mr+YXv7IZ3AphV9YDERUY0L/fcWzS3DC6vZ9IGViqGn9wyFtKGmBQu7BHo/b8zwxOoQwId
1fxMQHnJCncuwzCiiajtsfm/lZlVhDMeN6/E/MdfBofvOBNiqZdkKZE8FjabIw1nYKkecB88z+gw
BufFCD1LAlGqOITPDYUvZGduuU8ar4iC1oiNms23Ga0++OT6SQLrRJKJTFj2rkejPxCUd5Lf0F/D
aSUufI5DiRmARzNn28P7wXvkGsiOSIPqFdLjkMApC1Z/9K59bEF0QxH2SB1VJUkIO6NswNmZ3PRC
JJcZsnG7v/a+Hy5/Nxt1mT7WQVi+GtDRyKovG/sOZDdwn57hgNUPtCg9MGdquGsCJZau61+nzbxR
UYpT+oDFDpUVYvk1mO7b5Yv3UMw/Y/ExcpGGi9ZIg4jDutlaZj5+zBDBszunFaQ5IFiwoyREXHpG
O4sEIBPVzXjYsgU95D1+d2kIjik86cfUT8/zxs41Noj/ogghlpCqbrbum+0w83xXUIWIojyxxsHQ
ETvjR0kV5HvZI4LU2IScUVmCZnEriI/0Xp4QxuQP++PoqRkZxChfVKODyIEfrGLoD6vwyZh0MA2Q
iVE26pL6Ktvx/j2x13KJLZmu9SlcgAz+qhOZXuQ9e86oa3iv6RbJO/3bQWnQX5GJl/AB/bz2T9Ek
j134kqna0UR4dThTJcNPCvxdjcdJNRfuobsn+slPD1boJCMXWKh8E0xdTAO23/4BcB9JmYtkU4FU
IH7Gffzp1DO2sWEOuFrHj1VBSFgINzxMk+NqSI1hGfL5swtftnHiy3CF68i8t17y85TiA0iRwZ6j
rttGkFB2iwOLsWAAVmk0lHb1rzhhakKmBpW28kcYcgW6m4RScnv8nvy1o2uYyamszKfsXW+0pqEr
RGfEtQLqTgLutbFRKeUgHu6w+jaDgWWfZNYqbYREYZ8yj3ByXUm+ZLgpEbk/iLYn0VdcSxKrJEuL
Affgk9Nw+RzdXC/R2ycqNaqVePfoAWwP87t4yKry9VCbNrnd23vA6RpYterE15EuyzKB6YM3dn02
SqtQtPQDGg1f/PSoNYWQc3Fr7lFfsJmz4rwd3gwG3HAFQFfMhf1pv4CXxNQIFKwejQFhjjobRAbb
1Jocj7jnxEpptwXlYY6CQancHJGKa4A5UHHebAbBQQJKVazV+MKMSTvk2ZwW9Uw2vY+s2UN5y94n
HAq8RvTgYAUF071Fq4GZAegdFRjQ7MPuLERwC6YinqREbfuCx+szmgUURqiSZxJ4oLU58ybiRgrh
ofrcFvvzF5to1uA9wHaOw13OVhofRT+exSHovUAzpO+F8RTF8vM2wSImiy0m95rWwflxfbObaxgU
25beMGK+hYlrPcSj3kOW4KcWUoMbV3s4+oiNLPpGojz4eC9X1JCLs4F8iZu4G/ryfU+PfPyseBbU
oVfEZqCrDzTvgpZYSxCDgzepfh1KWoppZSXRvOz+BUaOv/h0R3FI+NCPb2sY0xL2R5yEuxms0Oxk
cbo57cxIfzGAKcEZ3cUXaWrdltwiPLIjtYjXOMuApxiCqe5ivKKvKlwWYYXfxp5q/itvaYON47Mc
mUynpgsBNN4iaSU+ddolOia+wiPIjStLz39naLximD6+8NYmdHLDWrUxJtbTeQWR3j4VUofogRtD
gQXNbecoKUiTkJ6rsaaHb4ZHY+WAj8NLzKhMy1axC5IYS4GTVGMbRIvvJ8CNvxt8jFYiKFyybi/B
AhdXwj8MULe1Zd/s9w036AXCLm80Z0Z4mSDIWVzt03BK5vDvxymxN10GV5VnIb8DomVCWa6wugYf
mdmoDpQzLHimiP+fbN4dt8GwYWj0zrSoofciLgzA2Z1mV4w+A7R7k3LeSBFbGk03QNDfJKiz6x0V
VpuEV9q1hj06ECDwpXdMSdR1FNHp78VxBOEDzs4e3qvZbZ9mio94hvu5EfWR4cJa0MUJansbkiGt
GjdtAztJjdSWCrHnT3d877W0d/ETn6MW7jxPMbW0E8GaIFDf+ZstrDnyV5s1DKu4DT5uN0REiaOu
wiljNSeY9h2HFaD17hyrlZqhX1Ox7Ipxge6CFv27NyMWKq2COoCCUZ+lRSYNzkwE7OcS/fMeyAto
100/puuz/9ZlQpKTfLHW6GPBaDZg/I+g1bePa8qDjQUyHBvWbsqD2QMkzcDH07D78sSzHObLmIIX
cKACGW0UaxCfETaJKNRmm0ySfd4rlaOS7deMmpCem1u86HPLflLxSo93z/VmqDaS1SFcM+7AQ7Z7
gkj4EsfVsRi3CmSr3Sxp4UB167nh2+1m9O1384/kcDlU52m8qZTXdkU7gFhySP5K+/Rm0f6/6Qt7
jVGccQ/PxoT9MDaie8UkH0jDCUuhuTJUhrzwoKrhCEaI5xzYKGuHLx6rxNoBa2J98vmUzdteYZtD
/ZttPvH9wikrXB2HicA4rhGzx0545np0F19KmAqjcKR7r8pH0mdPPKkpr59b36lDXmas5M5HpD79
/R/pSeAy6ZRLfoXO41D61/3VSCur3A17ndEaJRdp3jkIurHz1li1LV+vht7ZnFHGxaO2Rk5PAzMk
ti2v6ZZzp4gUj3/eH4x61gU8XhWw15taebK0t1Th/BmW3lfqcWucDd4tEP6dl/vwOw8Ma2zjLRyw
Pl0pBFaDRSQ7YmRtFwKLSwQAy1kwcrmKQKqeGKPVx4eh3F8hjmjKcZ7+BG/g3fBubdUNV/b5m/EX
ch+Iz234ej6btqRR8mdU6wzhOkadun5toWpyK9bhC3fxn90mswqqGqtdfujoZJ8FR8zHYY0nBnSd
0qzmhyGKdwE179Ui+P+aEaIRPISUFN3VofGDqVv7byD+rfTAwO0gNKXrBTbv+RNob2IVKpUjZZt6
maokCh0JttJBVnPKvLoD69iTyQJ4goMhuA/pozhljfGVGgQriyPW3eKnV36dpo5MdQFWeOjbfTtb
o1y9z+n1sISMiK9O8KTPDE6rcODTsbwjxu+hMYmujdwPHx3esJMQj9fLETW0L2nJg0iyxg3byv00
36snEev3HQQGt5c3EiBF/FM/jnfUIviwh9+4szGQ7D8k55nMG+E1deFRegusmYLJKXMhW1cHtFp/
tZg5vrNJ4FLJ/zCk+yctlTzf8rqjLX6n0pihzJ+qUv8J6h03GgavMq3B3A/E3aKuTRJH0NoFPgI/
VRAZ9CtWViEbRqdB/ClU7LG7P9d4kBKdb9MNH68hv4dWs8J/zwPKgEDpDRwHbIBOPUY/ofIlx2bu
M3egReKDjumpbSD7X3x/nf56yk7iQ/8VaM9fgGPIJjExFNi9IQBrpGJAbNWKAaoKzVkirjneCoxm
DMu+lBKkQrZnaZX4eH+MYTtACyAn/dil6ZFy2aXxuWaIzdaAiM8IMJYoxGk6dP8ASOAAz38DQeeG
MRpaIP06fik+yHAokvQrnYWzD2+B4J08NHAAHf3K9sfbnbJzJEsqrQiw4DlNTAp3mvp2CZS3+Ls/
339CQ20DxFrmuE6vXGBPmtWLYz6ENc68O5GwLG52SsvEt9aN6QoQ3WV/G3iSJDuobd5OWZYp3t5T
lJ8QGnbhPfzHZu3SsvykZ8Si06qXG1wJ7Qyy3z6u9D06dng9ssOHO5wBqHswKQyTKhc20NEItCFE
djEBSbgxPIrqG2phgAg9Xxs8DmmVIqtgd/gD69WISMPmfJJKOtId5ajS37CC6W5pq1JjLjQmYnen
zjXjfNO6RCw7fxWYqoEUYYb7vdC/lJOo4UkdB9Gsb5ya3tKtJ/x1FMqDAWWa1s0Ciy05ZVL1bm8Q
hKa5ZNN7CeWhEFxo2BhxvyiYrwICXcya+gpFAbfUbJ0Tr2SED24KKc4FNrRKtwL4Mc67qI2o/IfO
p+tP1CMBImWbq7mFYdBDOGAE9e0taYoYB3olVnMAE4T6Qotl9VMjhqfPs/0kIYUF+eEd9xqXwSox
qztn2QFP2VQwQIABbKK7GBwbYkzp9frr0Bc+2FLwPvjonfpLlGGQeUv5Pllpi0P+ogZdwEdKo1f3
Pk2EC47zjeu4Qx4tpEJ4vMGFkqIllKB8Q//mfJtIViHhiJTkMBOuZBoTDaYThUUbqVseqAb++i7r
75Ftk+uYlKFnQkU7UeqgjlFq0aXEYfTSATTyzQNo4nB92RkX4VScoFw0wPEIej0Uklzdelo7f83E
HP0sTr4YCck8M6e6+gPhaIGsAz+7cAkhpVaCOqWYDF9j5wsfS9QnlO6ThwICotbAcSjTJd5M/C6W
s5QRJlyaXoY/aRZZLCz5VUr/CH3cFikAGoJ5+LPLo7NQYrR1wGwguP8l8gTqryVHLl3PGoVUuhW4
jrjWtr71UC9ov5u6Wd0dfMqM4Z8KeJE4IR5cGWVJLZ4qsZ2vxRI+3wmHxF4bWUhWnO8MMYud9CQZ
VwVi9ETuC60dbhrxusDzWqY1DxT9mI5NWPbyBk/yXRVL3fuabSman8q4Yk40V2aCLdGCN5TZn2ve
xhuVzLYQbXEz4Scl4SaN/Eco++zc6U7CaOrR7zje6P5c3gB5+pDja8PtqolxZgdGO0gogSTqrJBq
mjAJNYMj77u0YUSPOaKf2GlRLtovz4bZEDEPsB50s5ofbrXrKNsr554+LcE7vgPplNvohhljjyZL
sl93Phk1ai/5VWD3wOWX8mt/7ag7IPBsVjLdEZcpi3DnmS7WM0l5WMVHRDBRFgpB7gZrAuvcuIJf
/W77nGYbpLDE4mXA3Y66cbenRs2MK998/Nbk6ge1H+w6Y/NMCAomh7yrmPYa7pu8cMubJHA2KfWz
sPCuCNFxQ5uIi2WyppjmoWfP+hKIUiUDtQ4AhCU8HSBkBSc+hwYz7KeXfo2t/8A1mYy/OBaW42WH
8wvyaUFSaCf/yK0bAfRkO6gQpYAtVbZ5cGfZS3/Nb0cnxjQ7/CiEZaW5fX6fk9auuPe05W+zvf+3
pMem+WRXabSoNoT/8sEX+2qZMNWMWAnEU99DB5tnEiQsOlh6FnNdd7J53vXx3AZZsuZDjq6HnfN2
aax/1+SdZbkDM8MEwKB1O+t7+naRujV+SNiDKb0VvZ1p0YThBrhrlTFsUU8uGEM5BDqWaWu4v4nw
cC5R+tDQW2dyGIQ7ixey2b1hDj6JJ22C73Ozh73dUI6lRFF/UPmeBHZ9MbK0MI9Rkt3ZUGv4QWLf
TVYVdj1mCt+71Z90klLc+rKebd/0eu8x1A0sKwwzvAzCOyUmQU+BsZRWZSDLrsyr3exiGPdySw/p
9J//UD7yDFVyL99g9Rnba1HwtxJ7LnksqNoTK0C7EquhOMu5IIdB1tDELRlGdug/wve7Oul20/oQ
Morx+/HmlPPiAtfTUe7bEc3+Vzvj7L//oyx2BMlwO9o2K8aLG10uZseYHRZliul6uI1GUBwBohVV
jvxKBvZNgXgOcxxswsoX7bmTXOzbnRdcNQKEYeF1PUTcf35RNMdTHZ0zrW+mdT9tcEPIwUvLTXI8
znelxuSK32o9GCM4xnopF602WQocTz11tfnyo+D2r6bQoy2hPcBdICo1SyI4GR1rLpjITDlZhEPv
CFBJU+zhk3LP/gCbHeI755rZCm/jF4giLKJ6xwIeKsbqUWlH2QDyQnOeM6qlAasWhFQyIKy/01OB
kCDOp18g9RAulQVsfGVKe1cNCzorf0a10tEu4g+D+pcUmcaQbVXFrrix/LQ6wH3V6xUHfktBv7No
p/o3e9gGOepJpLbE6c1NMBv4b4Kvjyanqda82AFsnWq06TSxy7aoebOIME4uG7VUcnwxgIPGkvwd
o4+ZF3Il0+crL0x4VGib79R+cBBH1H20H76M6oa5Tc+1m2ii83X0M0D+yqH5rwGwl0ADFPd05TVO
Pbuk5tGS04Da7VnyQCWENVuaqbCeODHGqRNJygB+m6msrGOL/wcbzbh1i6eJsgul8twG7kHhKI7+
ghxph40n55OIPohqZjPbnBHwCIYTAjsnwADFNWD1XmXuu7lBaJoiBmX1OlO9pTXygt8vUqd4kiMp
yl+8WAYtIjkldS0lYHa07Ag8iqMk64rUEVzrgfTSHFqC243grx1thdu3EnEpbQj7jfDlXciSxjmN
38Z4gg5PdxBnbNKlTckLyZutuM9OxoaGSwTPs1mOI+Iry9QpLygo0R05B+F4dPPuEoh9HlDDZN/4
cCK8UvG1YCSw17avFL+SranbF+7Eqaa/lREfb1X0qYRjg+g73X+KBjUcJAi5u/TrGkqRW9KKoZGO
k6kAsmcN74hij6GaBP6X4zGVRmj6yB/DPmrCiLG0TeTEpTrqQcMiHzqReaot2Knq8JZw5hZHu3Uq
Nhmk6XeJliezhmr4j3LCw0hbEYlv6LhOgmTtIc7O8UktGXEeam7zll1U0NATyr5mTzm0UETuISG3
cgit+LkppFLO02qjLUt3wxz6n8MhiLTzkWqS1dV1WtpVgsMP/FXXY/r78eNpbkd8f5Wn5F5FZUdR
1H1jy85zdZgzRIX9nK+DuV+RA57njvUqkzWIv9B84ZngI2WVm3qjVBnHouf/xQVQd6gDpsWRqEpN
pGa2UgpPOiDVa6T/vFAbBBoQzUMMb/V+/dD2Wl5ZKDlGYDKtkFc1jdz6gHfOP0+b60jdZKfzOdSM
ymAU1Fo8LlRLYVRareuImwqAXOdWYiIsjh1PkMRBSPujt40Ls2NGqpLVunu2UbEBNzJv03OiJDK6
oyrJpHVTilpjYfgS/Hr9mUNo6PLwNn0MB4ifbIc9U2aYghX2Tp/HueH4DJaKAwg8645lRBMSSUJE
3XeOUC9mnj19pJ8k5W1bT0atGdTajP/xuk6EbtPWE/k4gP5TS3NDuOBd4ikZ/XsCl1VTWiAHPjZ3
28MfplJOmOZWnYlrGdAOdS5YQRkegxrddTWMm1iYQoFwWNup1vqQhqXyrntuKeCAfNeA/ylFQmfx
016sXvN6kwMUjn3ZOw8GSD8NMSB7AsthoW3pytEf5d1dyRag4vw2gmOWdpS1yTRBSkFOrl5wEjYR
q0h2Fak+VjVugTPHykuAAoVzrd3wQsWATliYly56wYvZ+VrrSANVWIk5m0kFqIHPK8EXUzjiWsYC
Sflk5j2dII6NNi+CTd4cFj5nxJriLMYSjZYiEugUJt7y3/MgR/qmYoMJ97iILw5XAjRCN+WsdAmV
Kahzp3Zz4ug7hYmWE+/Hw1CEvkujnFzZERZOd5YZNepsKSNsKCLG9qGgmcnpsgI7yqLAG97AaLWA
5kImLcdeaZpUde9W0BgTgGADf0RL34cZ2oJV3xaSRklk1eR11d5lNqeXauMLYbAjf6qQyLBial9I
QJt8bU/sglnwqUbKHVUz7pSRvUcmDkM1VZu19cLH/TB6yarTgLjyTpDwB14PtNPOF8qVQ0IETMZp
DxMbQmobcsrRE/VW5on26eq3dfPbbHd2lq2W5f7TLV8XG71k2uF50YwE6UNuRndP+lyvmeLERxwI
lM2p0KEcbsoWbTqmtBnfoHtHeXfgFn4wbEwCatIteaZkZsmi35glXLwSRLWmy6YUhKGreDu/4Vn1
tiKycRnST0OB4q21ZGYDwoETBJzPg4/UWtHBOoCwwSkXGh/E69ruu4fRlzMP3xuo+gSJRxS5638K
ePRpvicnTZaFpZT8WhcFc8b3aRysMSCN+qDy25CQok37st4FURIdwyW/wy/1fqJzaIx2nVLDf3b3
0TavrkyHSFEwasFoVmTEdJVQU3HRSK8u/WcOmZXd2NDX7OW19rYjKFLTSE0/u/LcdUaSUd2nKn5l
9xtw3eKGCwd0gKDtmvTCrNrhoY6q52qPLC1nSJ8NnJ74r3FXCJOlyNYuf3xkh8tqXO1i8hHLTKrg
yW4clzDdWdvjKZlIHl/nRFw39W7BeMkp1tYFPJ6/PPOOC87Fcv5ge4KVvVypyHeYolNbTUODMZX8
zpajnShYtnUG0f7/vbZfHg+DOp/T+XBkOwD6yb8PKDD7rneyLO0mFLHr8i58L9mbY+fCyum8PON6
e6gXh4RNEtmEv2sEWIAcbxDuZCjQ2I7EQfltSjPmTpW/As1AmIoAz8czQTYUoCnG/RTTL/PpFZ+v
bz+AKROa3QW6hBYLuF0oA3SyUDQv7MeFVNs0yMmNSJzpE5t5QS5AiudRPULhGzAZ0XmG+kfGJpyb
Shbg5vbTixdCDJxEnBNbL78XDX++JPJJkpgl6Ux3/+lVy8JflFWzLDpkdysBlRs8n8NtgbD0rm9q
GbCYSNOMJFennh44E8lHhBay3yPyAg9wDfBbrOde6RuKfR6hnj7imDImlOXLwbfUSdV+rUf3fA0I
TC5rvpImNPi75scNu85Zq2Frji3uLhvJGVXtNkvzNj8ERK1t60OIylIZufxa+paQeZhiZwC5slbg
6R43ujpaPYnTV3kukNXdRKikymm4X3UpnwDexIh7iMAHROqcZ1R7XbShUlJT0MKpjZV7P2Fd7Zvj
jxZ18nJLDh0dp+PNex4HMxUAIgfAaN5/Vk8Q86VTnx1CK24IV7p0B6tsdrIeDoZuXF4e75u4JhSx
93FQRiJaguISZbFSPYEYFx7BZUM2Oj/AtJMY8mYPwFWrR+9f2RTpR71Y0IOcNh76ah+f/9Uc+XoE
SByCGsD47/kv5NI3Bv6JhYlHRCK/OYsthM1mvNjtuR6yD5T2cbAzsdfmxkomldrc9o7x4zZ9lTyD
wzjsYrpVbU+iOLFq6+ML1YfjlX9/HT/v0VlbuioEc4Jamr1V4rVihH7GL9bUrk9D0H82s94+AEf5
syg0hy/XUC8XJMIQjuS7lHi+IN6cprWyUk5YmXtnbOQ+TF+VzulYRoXGE5za3oZI+4AxkOm8v5NK
qgYZzLhxR4iloryVT5MMUBPf47vyJjnOotFDP48qNGrR0N+6Hui7Uu2ity8RvofPxROtkOACdAYq
jf2XDQSNKSkT8MNIB9ko4DByF+t4tJYqXHiEPvh7egNlrLaa5XvmcAhA0P8bLeqph+D0i8OMUZAe
8EZQS60omWWApeh8rPyJHWzmwDij1ZCM7iIdA3Chr0oO0NlpUXX3kjvO43inPZnqeXO1AjSLhiko
FCfnD48XYvmwZIns+ImRauWPJ+rNOAHRrX/ARPczJ3W1hhSc6qH3ZPxdmrBM1kuIqJTUNd4avGmg
Qwq2YaNwxBPDDzCwrHfhJ7OKuxdr8Q6lRp9CvIruTF246p9smgxIJJwx8zSWR2VK0YjGeRsIJ+fY
TCFsZtLoEoYFGjYhwE+xhmhy2XYewmBhNC39OWvcHF2U5C3axfd+M1G58ZIZ5cxuH1SN+68TV1P5
6CbP9oUTcLYrpINb1zMTrX9stTM56CArymqt69bsjfi4J6twTv5SXXQ3ol5aiNhfUqzzwO48Yz4J
jSWgceCSQF4V/t/pMmaO8tlfncQmAtUO2RGEQgQv4+v/NmrOowO8reKhXzRwft/sZa7XihQot0ar
XvhJRevV+2KBGb+qHJc8pBXTaMXX44yxAN8YySYJm2RecIpwRrras0c8RIv8r8VpHFWL1zUJjWUW
qRG0T9mghfv7LavniiheAe1P0yeuhCx6sNxjlbv2ldMN778ZQWMwNcs7H3h2bBCsapSUMBZu9rr6
8rvCkA1xGRPFxMymmBROkbqmYvuzIdndjTOM9SmkwzQSqvESu4Ni7lj++jjkbavQy+F1wHzpmD4I
7d1kzy/QS0TP1RwEmD7DXUD9xl6VzV6XmCRtT1lUejvnxEvQt+55rHTadDH1y2nTPx25QGuMVzWi
Eau1MEsm5PcddYoABWT3+tlegXgeW6TtG+dwDzAPuqivg7tx44P6FVTS8WQfsYAYfoHz9gVFTUcY
NG3N7iKQvIVmPSFuB5gSvKjmWwzcQ/jolqEGTBjdLRr6z1O+z4M1V3Q9LZuUIXiVpStGbkmtRH8O
b8mqQxCaOyA+iyRqOkx56Rq2kEe5d2/Xxzie+MSjPpXbezXlXsiqG/KOid2aiYkVpXrlLRUpsxDp
jGmkHgD4W9KZol/heXmdKOJtfIMiFRXNSu72cjW11YePiuyTzpMb04ceu8m9oHgMDV8f+T0uQRJG
ejbZxTzECBRZtBjtKmbnKEzITTZMglEXoNYJXXkZ+4ZChiKgUk3ECTguZauHQb+7dLjzK2fBQojE
dCIsV67Z9QnFRB56tm0Ftdtnh8g25bey5bzGB5zkqoQJaO+of5Tq+6l7PmUpJ4jhBQ8nXRW8w3nT
ACnDtrWFAA3iJeJS07+A79rjjxmA9v19Ws9amKlOBKG534xCFMG5p4y4qyr7TUaodFT83rQM4p+n
m1EUiUVT0SXvndt1jb8HbV0h7fEcttR04ENlqwIUv3rd/g1u50MGqjfDPlsu6YiW3tIGHxKI0AtG
d/woMWmJbdrVyTyFy0tuBhN4AwfCtCm/FmUdXQt59zxTjZ9He8EZDeZFKXUtkRwP/Z1mDh+XNTVw
00q9AnVi435ltXCrEMWfYmkMgfDPyM4otVHAZiyXs0HhWfkRt9XoQcbrRyQkeWy7kfdQXAu3iIgF
VFaDsb5m0V1ZrYO4Qy5o0x2dBhB2d+C2nvaprYJPQTzGLLf1+H3Wxmygf85sMEggBN5gCpWprlct
ibRjM8dZjY/PGEB7gC7j71m8TI3SVLCAuKQMyiuEQmjOxydRnoxuoRwHYbiRkcXzMnFrdJWsbrIa
eYD2zj7FhhFEE9cGcfb6W87akA2cFs1zpbc9c/4TZPHs9dSA3qAqb4DxI3GwFuRq0vasuPuz+fx9
JGZUCYKhnfJN0N6vvpbd5QXKnLXeWeNTr87++kLLXPdG6ABe23dNEAYJqXBBLmVicnZD5SC1it/4
HY12L7IWVjEeEKXTsmOVHIolZdmCnBvIXtF3PpWhFTM6WXBSyLTlugks2jJnYbHJZAYp7LHJTqBG
ppLo+CrmLlElayJm1ixR0q4a6bIXcBhVFzx8/VTvrAnPbwQZNEnDR3XvU6Rfetj81JR/fwwDkgFd
6awN0dZQ8r/VgTTKXvX1wB1zhzkWoR+ml2hxhapi9AZsywTiWtyb8Rby14jUAUtwybAGvEtHvSil
M0D8GwxTH8Y4OH4b3Mjb2vLLHnv0rwEOGiJXtSNADEbDDsOes9XIfuNGXXgM0bsCJD0vsRgnqdsp
WNU0MA5XYSqJ2oCOabAOKt0dtIDTo8EB2LRO7pf3Rrx8XXCfP3mmAHTYQo/1DVzTHke8zHCgXFK5
OjTyN97dw+EXVxidQseKcdNM1yZi5yLuYPq4SveDJCdi+4BWkVGHiigFvJEnXN+DJHZtici3atCF
hbfMgN7BUYs+Klz9ZMgtxlyxKzR8z+uUUqWXn2y1JylvTNsH6jIR6L8+thiiAsx15i8wlSMUXL2g
Uo29avlMt4J5hfs7YLmQ4nhMU9oyivi/GoPdjNhNmLKUGdCA6qK8k/q8zUwQWO02veoMfK5oZcOL
/xxt87JBq/c7wBuRZawFm1+SvNM2Ym0Ml7etMWDaBTY5+GicSHI+/wNOdkRJysFSzo/g9lSjj4Wc
OlvUeRxoq6336W+0BeP1Nbm3JC4ts6YZ7NzAqTCAaHPhuPEvnxSTRtrxrpgv6RnR5+BfCfzyRrCP
+JUwxXeV44MvInMf8Vv2zWPZJrJtynm50WtEtnvZvTH+56fYwgiyq1gr2MgBLH4jtWIxE3w6zdGM
SA+dYpGCV+aQWHltXgHBIc5KcaXGUSvxRe2NYhSdbALJxU9SQeICGOnkvQxlXNqwct64b4mSN/BY
E7h+SHkjI8XwjvB27k6I+WZA3Ty9SFoncUZmpTilqEH3uDaFEz4RfddlsCJW8yeczlg4A/CZVkUj
8JZwo34qo6lap1JQTAR9l3UJqo77DOL4xmzA1oPjk+o7D5VSNn1dbNdJ+K6nqMiT6LPsA0igaKXA
Oids5zrquJhfxACF/XUcTOCHieLlJ7T6+FyxCz0pWTxyoHboG31SpTyAy9gdwExoxyr+Js97lDXH
gG1exYtvzwpPN+AGhQfpTzL2WAknKctFkm8raZqcxKExlbfAjDTteIxa3IJN/k7M1X75i67T+fJM
Z0TH4ZePQR7+WfWCaFoiIajJdCvBFbKeshh7mX4JczsjinmYMtz5C9tm3iVcXnTrgXGSQ9emYH8A
xMJ00d8cAhe2z56Z0IajTpC754ndnkotd7GlG+PX6uwlwFCM+HZjJu0/ZfDn6T9MfarA5Dt/XDj6
ISgVbuYFTvPF269UhTxqpdbyviOENa53M7xRundpfzdZLwevkM8jbZ4UJvdM191zw2hWvwNetoam
Z4tYzSL4apn8B7UfH2LfeKe8J3wqnW526n3MmRXnlL7J3tSHXjgKjDXtfa3OGozOUGOweBCoSo7x
q8SINkUcVWF8mW1W6TO1VDDJS/aYSHB1Kxk/Nf88ZsImY6rCRvnRjvzlfg/wXHC07W+ZBI+Bs8G8
8JiTHjBOYlP3RHbAL6nPMVsJ40lH1h7VK/b1xg93Erl3rwVkz9U060PT/PHJACuLJtQx/d5+dx23
bZlNyMRZ0SL0EMZKAsj6n7Ugr4uMvxDajt2URdzZ28FXaaG4zPZSM7frnIbQVObWmMeTUmLnhNZQ
RFZ1iIg8i74nP47FPDgN61XheUeYDnLBGPcSE/EJ3Z9IpOMdeRdZhYjNPdCkETaFVcsW08zGhkkI
YH4lJ1XPpmu5lTOvL8TYKywITvympDULG4UuKM+eKc1ukTAymiuDs1D5XrEocVEyVblv4cLT95XK
F9Gd+hbUcLOKVQbgJHuhEqZVZn4U4R1gFfkb+qjmwD8YwKfdqGdG/BCy7QqdLPvbsQov/z5cjn9R
A+7tYSaoguH4HLsASrrawBAZ7nYkgcVwnaSlFMQ0PdGmQrd4CL6iDHNvsGJ3Sw8Koe4nXS+xwsyG
MTVyaMkrjubo7EzwRJ0/wMSZTzpVSWXS3N+bYOMKiP6w1eTmy7Id4dcwGGG+8l1UX5fWN1owR1a3
AfoXJlNfw1QEqJN4ole0Xe0Q2XleRnMk4nvys25ctvW4UvIH4mhl4lcFRitcPOHm7tvNOG74NCM6
L0DSs2eYxxIchEVe0hv/rJOewonE8M5Opl4/IoSUyFRu56+H/3ucBpM+Mi1dLnpfbCpr8W2Qjisl
QeUrfJtAEXGVlLUfNG/gfoGIubHonxbYD/EWWeLDr0+H3wSocvDxHZAKuEXn7YD7cuNfDBd6SxrD
jv3e+utkoM0/6vc//aq0AtX3e26UZ6hxfZCo6jXpVqeWxD8Uj2F/MSz6dZuyZHk2YtPPA481Vv4i
K9n4XO/Dz0UXzmQmz8iAcgPdeg3nZwnBwfvmH3TWSmq/7qOAZ7gxoCVt0PNNzCV5jHhFQqM2flbw
jH24npXyoE2dTRveKrgrd2t3F2dklf9imM97GxPIR6bSYaqDwEtiW9/i+q0u2FjvuAdgmJ93V22O
aokk2BGH81jKVKOM+FZuCoqz8c5fVtGZJO8uIgdjvo2ZSXOYiaTwjYiDsQHYl2xI1CKZT/h0KDU1
Z5895uToP/yEz6nWLEea0x24fnwI4WOjj8FFgBx4CMhBWUPWgGewRb4gCReTAG7IsBN4XTwXDJUt
NQS/VVdHo1gCGT9YNyzboBe3NonQIKItlRXX04bPkzLItJyDY0FlFzN0KbZIbv14Um9tclH490OR
Ua/qYY5v2wnt7BjdxYpAPTqOZYDTA+I4YU/S8DLe6N2JVkr1HSqVEd8DiAUUs5BQxJII4Rxq5O3p
e6DMutBK9jhxQbvLHBb2wj32VS4+X44j4isoa3U4U1tZYZ7rTfaW8LRLRPzaTFut911ugCPxtQDN
145EK50ivaQAUYcv3CU8VA2fB9u+ydJTXiimVOtVvDyRkFT43BQBQBZiZnSFFrrWqJCnHHxirGwY
FqhuIZTTVMuni+FpKawt0GHb8foO2dFVIIQrvkmrxIkVrf3RT6IEW1/I8j6IXTOPc8HaFDgJv8jt
+Y5klc+WxeCZTvnmNPHZIWopGuGz80arKeJBUVKtf1DPOKhzAHKzzMPbSO/yY2Cy9KnTkplwEqo6
OA5IH56UOe1sVfcFNfua32uAmhZOgo9wcAQ3lVnnBq5Ta8BPOtK6ejHaFi0cyeOLH+hL4bRcLtil
YCx6FhhN2XxjxhkVsargvv23suoaz66dGAVfGjagP9vqg9I9241Wb6Y4qtbTelsPs9PfTUeL7vgI
NGFc4to6COGCETy45KGXYqTWSQkJyAsaeK9XOPBT7xGN3VNvLcdBUCmXFWltr+z25BdxG1cfAg0+
q/f3iIqgdVkvsbZlCPTjic8rUH/zEATfsLFxVAhwk+Mj5eU21TWOoy36kdP1dZpeWDZotaayaqrK
nyTU8HWxne9oaVnEEFCrS7MH0sxuyz6p1kJZe384Mfx9nsz8ETSo7D+l5mqZnR0RkCW07aIG+qig
yKXLVLg4MwLw7peVVAT25EZnvHjQnqYFepRIaNwMlzUYlBclpHKqssHfbI8b/cb/FqRuLyI912OO
rjOk2lEPbY5WQv/HOMWXSA1RZhsRH+uQtJlOuceyZw5ZyJAD6DX96KWXe1hWnF9ucd7+GsGfDmAf
5Z+1QK0ZqjKLZsEBfERUyHZid5Lsn7waFTPQfmVUBDc7X1wZ7jV9lwMS/tL5ZnNivxWaTacQV6mW
I27xx5i0NEOeDnnewWh8FZYFdvmabkKdU2OjA9MjebCeQe2O+uDcps8eqYI2pJ8s0iuXUZ3X87Sf
NfqzkiCQm+LB/cvkSAASsY1qSEWj4jqjcEWiXuZuSwdNxlXWCUulSDFOFyhwdW+Pcv3iQ8zxcBBX
YzKCQ/UmVlUMFI5wZmK6wKnHke7YKrCTEPCob/vcxHq5e1o9oKvazF8eC1KFBe+C5R+cOweQxD7I
V4K8LlMdIAlh8m8ts6gOSHBMGbugv0siFJNceAD9kwCMjLkZ4UUz2xB5wj+8AoMwd+FH/GVIp60R
xIzqi3TTVZwUVcfKctKN/pMOaPIB712QqZlkUwcHpfwl0YlLmWeguidQGJuNZGytpBiBKQ9fNZca
1T4/0s1kYyG4wReh9mdSMd1mzjMDC2E3FsGv9jb8g+f0wzTpGQXuXk1JZC5S7JIltIXuRL6IL7qz
R3AIUSFwRT9nlFl1B8LDHF+UE7Y8cUbwTTcekN0Y5Oqvc0NNDds963flnS7zHCVnDSe4bn3u9Wd7
Gx/QaS/8+NHlqgKOClH1pAcZC1c1j0FwEEDdwZYhEUX7uqx6xzUv3pq/ro18FICLJwm9u+wZGvqG
mthCShHKWZzvmgVTKQUaRJYaWJh94XdYl8LfmfhX0iV0Yw+Vxs9xHzqGwgzUqG4vNfjImuUtu8CI
fGEknou4LSZGSdgtvtlrm0+PgYq5AZ0k/SARJl0ErJvfwPokkNBvgtfJ4Z/OrwOpBXwqVPvP3vDz
hEq3h6ATjMJihpIygcUpP3Wui2++hHuHhnWdzzttvJ3HvsfSn7/EuFnh0Kqj4lYyD4G898Fw2USi
4nRXTpG4JCqlq4NXDTlUYyY+tF4cSLUa0lW62bx/ce5gL9BlJeZeUyXcQs1gu4WIlJHO2nwzoF6r
qllC2iwkuVvpayigVq094hyzGPPv9SvOsvZIlpoNoGLTjlDKjgQ4pmO93/cS/YFXplK0LNx1vLh8
BKXfax1x82OtqpcA6aO+BE0UBW3bur+bUz7vNXbrEsCJTsQYpIW/n9BG4vAYiF1rae6lPN9an5Z8
VXv8iGBTpLy+hgRvCNlh3ccHbYmadeDRqzqQ2lm/RE1UILsN7jiX35obc3aDME0IodWzvKJvZQe1
1SJ6Ji6UIDthYJ2ktcP44fQjJ8W51YujGSlQzcCu8sf8iEG9MRkX1WwihoGhD6KwVt/kuIF0Kj2q
bQqAm0WgILO0LGJ9yGMMzZ0SD+7oUudbhlfbMDwKu3WZRgwSqIoSvrW+fsKPV4Y27uuwfWaZJM1P
+MMPp++jetXRj2oM4mvpa7oUORSKUB/N10IGUCSeSVe8ZBOUbutd7TbgsRNqD6ABJFthHJ6Q1DO1
UaYhEqUhZ6fT5c9Y/7+HsahzpsIWlF2O7/CS6h6uMgjL8i0uO/y90ExXxbvtsig16+Msz9ydraHn
JcHCz8FTDtNwWQ1TZxpCqo7ywGRYOKVuBwsJiSS8j0ga6jN44Wte+D3D8zttPq7VuHwdtf+OKs+k
hbkO8BGtt0LnLYRE3KMU/vwEqvY4fcI0OPoXEHthmNqcP/qeAgrr8LYNT9ZnU35vR/ZOcTMafAYm
wc7ZL3IAq/jBGssHMRi//SEkqcBvaWspCl6v9vcEjjeA2TEYN2BSupfh8nyOnbBvou3fwCi4DGTP
+3MJXxVc8eNWs2c8SvdvpboQXJaZrD+SIeTkt3HJjvPkF40vvN5571fkvH32pzj2xYB3SoGNzelA
0sPRNMQYR/kCSDjrFNc7PateagR+4iNlsHDYxBVYoL9NTsv1tZ1pFC7V0uP+/c0bdFACdrT02u4g
2ttgWWHQ8RFFxtanwiIYx4bUsQdwoabVXMrUdo9FiNGjJysdAyX/wGjsocMndSuCdgozNhOI2Xp2
RQ5smUnlDc4FdgNOtcWBhXT6QM2qmYXJBQch3SSiPk6R1Gov7Nzz7/w7fZVXIWuxY5aCQL7XeqYN
UM6KRa4i6X4AxOoYgG7NLgvPALQTStJUiHt7aEk7cOE6Go5UU55x7oto2hQ47CEH5tLzHHdle+Js
P0919IA322mPsjJsfsXQcchREUdhT60yDYB6zurlF+bHZovpOtkhtwz8BXu2aFBpjxryZDB66uVm
hcdO3J5S7+SaPSSdVEX/l9FqlRky/oSpqG8aIy8d2MSr286HIni4ceiBBQO6KNZHWJU3E/qrRiig
K/f/ulIGxpHUw5EULNsZMdRWFQOfaFJ28XRmCAzVEO3RIKQbcMyl6DZ4fZNQOz35+6ho02rgqIqP
+MuDyIhj/rc1oXQwbm8h/CHxpWkJbRD2CSHWVc2VijJbWPzbkWLWbbDyrpUWxlGOZ36xdpHMsHx+
EhzN8xtc7SAwj15Z5mRZLaFmedQcGfQGsxfY6l3sJyWJzVAb5YOGcXPZkdHlgDmNui6ydSlWNUSO
SM0g1gG8z3UypRM4qjOfyzE5JrfsSIkjXiQvg7suDuCCwDMSZpKy3NFVdqUd0uKKXTbeBAycRYWE
htwA54ZQCQnm6SuTLhnmt3lzNghi4Q1kECRXhuj7HITmlNgoffxDD/6eTvHt7A7K7ESHiaxXHuHL
9uuwcaaO9HlXN8rsF8XbUM6vhs3KP+T1veaj23bCHQf/dClliGdo4OoI49ME8U5aWCUqjrYqbU7O
YN+YZ5e5TqfKGpcDrxzbDARudHTDHmn+JQP2y0u4OjbSDyLcp1exJ21x+bLIWmt6Gjx9OBAuVAVo
oVQGOfcZAC1wH8dFXJd/p/FH4lENnF27zZmHjixzHLXFokhIGBa9VkM/ojWovOjZR07pR3EHRJS0
wDKrHkwWYrmIQIU025alFASDDec6zBXRCVKQXqyZAAKOcqVFWbl2g3oC0RaeRfBWUdfdl3qhdj0Z
WxiX0qc/4gsEXqIvgVhpws5YySTXUpF2WQCznV6VN0obDvPMwqOBlpeAAyODUR8vqlNA/jekfQy/
w2u0VKSpkH0/CWjrm03p+R8/pZROKJYqW31zD8hfsCjwQLwwPPLKzhmgcIB2NFtt2/KY6DQMRREf
/YC9+dAYSsrELNo9+uzTBbIJTGfGzLdFdLtPUaxb7p95jPgf3ZvHR52EBiX+9Nag1LcmNrJ4NMf0
BXbfB/cTPK1ufacFZQAcOvJZ23JzJg2j4/yc7gNw+i2lbAvLcm9ITafn2j+rlG0jBW40I3Fp6dw4
mfDJw4GbD4ZaghcC3eoiCSxkjjpFkoN5J0Jk3xgidskwffeyd29f68nrSa+2acWnBd7RX+TajB4n
N2KhmHI8300qDt+NfBVOekw2ej7bOp0QHycC7xt5Gg7H+eseI83l8DKDgFqjmWTbOTFN6y6PxXW9
WcjvodqzSmpfa1R9mBMjjyXYdGmMwaG9oTwTakzd2HZynM9+macfTTk8HJTnag+GEH3EDhknwH9W
S3JwXDw00rP3PeZtcdVJK/cFp6UH/yfLL7+2Ml8SkUvk+3pXHH+dB9BlUz5zCIDRS+q/oV8gnMvr
4usWdagWs6obFnczhKhjcllxXYEVBOofULSiqHETTWuwJtpFAmbkRPRaFngw+EQAFPHycSOfXIJy
CEhmg2Il4dDomgl0ekeOrDgXDKab/kSMFw4P5ZyRn6g22DbnH2d7wJasvaebdu44TyqhI4F+6E+Y
GJWqXfS1MEIk29zfvpj08gst4U84zNjGxNhE3fCVn2C3WcMI3TpQWxsoOsnte1vq9+53prFbqVSf
4Ns+i+nJnCPVeyTxNWWfoHxFfa5Qub+ObO2SLBtET5NCAwEf9wBjsBuf+D9m1gQ7BhrlQ8MkEZw7
hg9B8DCogey4HIM8UKqKkEJdGaJV64n1IC50Ru101Q36+vD7MdahhCLhDWEHm6q+UCi3JXM9kmMt
BiIgWFXiDQJG7GNLOgGzkNXpKAXGHDkGddybCpAUPPbmylJoR3XVp3HL3uTS3XvKbe9Ok+CQs0iM
XSNQqlK3E4zgWgAXIOd6CL3VQ22JhnOtI/+y1Geuut1n3QGoJvWFUO336RSaiLwbR6JQ4lUbxHIq
RXfZc70VlkqHXYlYKmYkfZcM6hCaqqJO7BilfK4yPaRU+GzH8WiXQSqDkH2zjwOpNlMWlhz5de/R
oiVW6RIRMsf4O99GX0TqQEqIOjCI9pdilpjDo/pybyjFzWGZqMAMOTcXyTxEp0BzvVW4pVegRpQz
TGFdHQzL5DuVMEvGCvbalyuoHrVIoUt1oUBubvxomWRGAhEr/JWiUzxhKLnIshHE6LUGF5qn8Dvp
6VFK5/uBbi9cT6EtHSUhO2bEDb1JTD3iQwATc0b+RSS6uSNOTD/YgSsQyWk6+9tROPnK/FZ0Dc7l
xUhLINNZnfrAHImdMM5jN/1GMamiK7YnaWYh6EC3zLXls+GEwe5hH+T+Je4FaK+saz6a18eRBU7g
mBRZZqHCPcl/Nc+54gr1MMLzeqyk754j/yCtfXvmnBbvUrusKpP4fnATquZqWV3nlpJaGrr4MI1g
YoBClRv+fQx/8gQ77KYapAiddHvtho1vaZmgj65ISnr0uX9Pqk1djtd2jgZzJpiN/v0qSEqa21O6
3MDmG7XQ/bupvRJTJwwdfwAsY6cAw6yg68ti3RjiaCBtsbfAiKP5Z+hYfgmFlBNvwm4at70T4qyU
N04iCEPNVEt8pwNRANOoY+oYEVgY3CMK4YSRINhvajvetaSvu4afzA1KSDvmtN+akyPFcmG9AFRG
zyHe1QeGRn7LeOMlrZ7Z/XFFTVm6MmiYSE+9rx8G4nqdFcRTgZiBeSpj5iLsf3ePZuQ7bYXPcGnl
Zlj4otiiVVV4A2/u/pbchv3dLue0NYy6cCYywhluDL1erBwkpCC81WhfSm0y1bs1gQA9GdsCJrOb
uwigaLPrEzwEF3foFW9HpF0tLmKPruKE3LdA9k4DYN6aAfmrUXk9tA9pid9EpSSdYnkDBchaupO2
63Q1TWugXn6bLZU09Rj3HIgyPU1+97jP2Mg350AfClthoeHCBxd0dlqDJTbS8/cfqJVcfsstReIN
M5FjvS/otUnNCDsZmaYM42bZvh8AH9HE5p89xvA+WSrDc85k8JcbDPS48Czmiqw/0K9KPKNv2Kri
vurNMdAgVJ0E/DwBZCZ+04dSGRElqaanK755zy7qLLE06DDLHiYPertVOIC7UWebF5LE/jf8biU4
XmsC8YtWdDvijl5gKWUo7LKRn5xegUbsjzald36UJcHzdJmIfsvL7OeVcT4zj2jkUw6pLD1FsbTE
D9YFbv6XmMnYNOZWX8M3v5/KJfpaIFKWXjuvfiCwQxCCC7U+hJCqC5rPjn40RglvvzXCM6wvJxLQ
X1Ez33OmR+7Bv3v3eW8mAZQTLTLMikhu2FBa2QL0acAj+4vIp8rjMVOnEmZ6KswwAkqpNNW31/UD
KoBAa9hV1zMsSWmlquN85piEJIInatLLtfR3pOZjvI46pt7TNbPeCcf5DPydQA2IcDrbUNAvMfVX
/BLb9uHIWlm8JNjIrOmLkVpoYWajBFpNPMEFiv3y2GkXQTiV0sBxrkUlN2Bk0uAYuj0QO5odyH2D
cWonE7jGvfziiPCdp6YojnPDYutpW7RHJlOcg+SXT9YoO9TacLwh+m+ChEX0p1JwvJzkJTJCxR9C
RTkF4aa49LQqucAfWKmgOkI7WN70b3aDX4d7yjaT7HvO3bjqBzZtu8carDMHaGJyIBKLdsyTF5RI
Vi3ZpMnn4ozzCy2zNkO85ytTuBWOs01CNzW8RyogE4kmgafyt3uVNHoFhTTNQIzfg+eMsbZ1H2qE
0GKtNMvlBvmhFiuoc1Vuuki7YsXE21AtswNZ3KXSc7qt7ay+tdOkFxtrzoMxM/yZ+p6P39AQfqq1
4ivDt8UC8tVbFlHf8xpF/9hqswlJQoRBHBcMvukq7wDN5OWhrDqjkLhMyPcJDJ1vY1P53P97jMdp
olJ9SbUWVtrLji+cegvb8KmF4GVZfAGhiR1lMF/xgHmn1Bt4XxLX0Faayh8ThImysOekMEhkHE0s
b31RJsGlOpoywJj6/2UCMY97KB9P2nKSmCQ18pT0R8eIgdP7vEpWUrw9Ws1iINkI6XxoAEdlvbkg
Wqe+AfnWrHPnlGsjHuL7U8TJWLuo/nkMO3kvOcgd/ui8rLnclUKuB05toZCPy8HR/XUXhta/YAk8
TOKE4mX0ulRcMb61y8vZHtvTO0dD0qhX3l1OQYZswNwP/zdU3m8rAqktvn2V5x3a/Al863Zw6sPr
y+Lns8aldN6QdcmVHpk9jyuNcD5YWZlMX+BomUqmZVtdEkjxaTxgpPt7crOSN5aawrgPjGkmUT/r
FfjNd1ulxDIFpzWZA0le2uAik0BVZcn+C3Wi5I+qthUmv725sii+MZyUuLvxA+HpRapXfrUJQ4I/
idJ9j14ngPSIYPzXJW8nfZ6qSXfA/97t3t2nTDHNMEjRecSBGeHtXZ4pk18L7M01ZSQHQyOvzeG0
XrmmP8ZspeXHIFoldU3zzYKNEPZWh5c7RCIyLzC1Gd3dKh9VZV2iJjMEoLPdShIocr1cyI13ukTJ
GGdg0cYYByh1l259h8AwQw0VoMxSOOwghnqxL/ImMEhwBekPNDc2fjLmGza36SlJjLOLMzNfZEQh
N3XzfZ1/vr6+wr5Ae6MhfQ+mgaiHoSupuW0xrhaomDeUCFWmVfrZ5aFOXuNDvx4z1EUmKQ3CnPW+
BZ/7baLoSXx3+Fyf6PZr8s1QbuNkYZ1hUQXVNDMlPHvCMzLOE38Ads89o0tv0if+qS++CFdCZiAI
qMp3y3PGmF6HYjHkOrc+QWmCGBc38jL0vklhytaAlWW70/ByJPlcW24TjRwWjfuk9j8oKV38TVDL
FElHPNWnkJpVwMcVtvjyzUrA3Mnj3N5vHEExpYpqOO2+biMU3pxnd1tmq7jgNGfhyXGMgkjxqjTO
ueYAJOOlS4a0CAa6YX5DzQOiD7MnloZ39r8Q6tPSneFi+lyNo1yJ7e4Vw14Ut1KxzUuwLUgQhuvI
6Os6V8dD44EMKl5HeGWk63tsHMXR/gZTS25B17t9gMOdJxVw26l/fMT+7kyVyD1z3EPvI5a4/PqJ
uZYTzOJWzTDZRVLu2iu2NJvj16NGyjY2nR/9Zaeg/m+fSqWPrccKEMzdsqjNRXLn2oV/1VWFmegF
DhL0FwSVhDi+EKoT3XJQFpvH5TLTKhrrSRBxogCjY0XNjVDBKGNc6dOsJWcfZPvSmCbOwXX4aNqI
zWlIYkOzayG/0lxZy3n1u8Ar+2gGxEFV+lU/Brmj3Fr422mACmo7TmZQaB+vSSsX6scrUwBiKA37
O0dzdjiecd0iGrGLCcpZ2sYiDKNcEFK+qoApi8hf69Az6LNHCP59Oh+I4Tdwlb8SQo6GrSxBKTP3
AkbM0+dfH5sx6rIXmW0tIyJPxdnybKuELwpqEEg7dBCJfFex27MdU3hFA8Mus/EsPQuaGRUjsc7C
pX9WMnpLjdTSy5GIwr1R+WaT8LZKhZyjjAeQfd94IyAN1DfiZ0IGx/HTFUxWQnyx1an/4lnSEOV+
duG2Up9uh07Pq1nuNFvx6qBSP3vXWs7kM9YllNw68z8tIxtwrwRcGwHNrJcENjssjHh1wFpjjvAR
C+N/VmqcDpwZfRtqcpse7mTFDM1UNH/vJunVNs3mDh2JBHpBaykoGoxhcc67vZNxe+U2khfiEDol
VyQxsAmCN8KtqSGeYtb3jrQtG0F1HFW6C5xmbP+8vhb5fqUdA9BjZOz1vcehkWJOA0JnnaM5sPka
GrIauZnhShhGFaAJl3ml+RuhWWpLhm1nK43HHwN5nl2QVdHMmK7YyVrTbtqL74LzHIvJEdT2wnSt
iyQOIaa8XFkcgbbnypjunh9JU0TuUCaM1shVjVOSYZZW2JC3cjbwfbg1xUXL7eZLOY9JBjc8mRdy
ZQLM7OuP5OK1Hoiq3tsz/n4V+rTuTbmdZcMilQNzj4jYc8MpZlJ9CjclyeMtTV1nT3CbLrNve1IM
wIG+p3ioTcDkolXAWZSo6T2klVVbzOklHzM18oE+hBTYzoyaNoHUPQklQhT9rksSyVDGZjq1W8+O
SI71TXqzku+2fQLYYxlPDK0Wv2MQ1vwvpbFp+oUNCJZIW6E6TbM9s3ykjSOfBebwXJ/9RqHKQo5V
mnS5MqW6aKxwWc0SGOnVmpjVW3bLHA/JzaYI6hy7b34u6V1cM4h3pyCMPGha6DvfIQGEsUbmz7FA
ExPQpnKdFhrmo9ctT8xZ6bhsH2Vmrxbg5xn/Ri5StoKhj3w9GIk8W+yZu3JU1gNAahNEhyEzgTuv
t5z8At34RyrkWeylNo1olzo6+8IPbqe2682siv4Ya/ePBtiLHGJfEZd+f0vpY2+SiWnVcowF9Mz9
uO6DM1BXUntZwLzoNvZqakRygQ+wItTewxSBoVpcbgXUY3enhs8HXIsb1Y1KUVqYEI+Dsa9BOQ6N
U8ySMcDLIvnJv83Lau3doUDl+dpofCWBEO5AzQt9s/wZW+xE5Vue5GmJ3PG6g2FPeV1ySaSKK+fB
y1JD+Qam5L3iA0wPRZoZ3x4aSgX61N5O5Hr+22t4hdBsWjbN1jNG7l/hzedIcG/tabNA8VQ/4WZA
ps797S1IevOAQxTCmtY4afQH1CvWA9j3TWF5OUNb6xOcIcssZqfgTZHMgBJpCojP7/AgK4W/f7a1
q6Yfxp1nvmsN+yY8jAoRxm6ieGzX8XjZbjolZ0mwncLmct4Ifg9jq4NzYl7AbaQVldckWQBY1HhQ
0fvFrFWKmwCozeLYranQU6q/PCk7HfLHxiOyoACn8oVmSeIeXymtHzfjK5mGlXUXutKe9O7jmj8S
+fYWL9DtnU0a5CPPFKKG/LSyob0oNDQDWejawqGiL8Bs5V1Cm7p88jm9SU5ZPorT4xx6oTx3aiHn
/QBheIVFX0GdY1jexXd2iYIVByw3hxgvRppRU5FPDB4hDqnedohqIFLq9X8WtS/3BTCtA17pMO9L
LzXGmhZnEnLoeHkaR2pbxBYL/ldjsSAnBlztN1kAZLaVVG78CxeLtpIOK9EqWkhiPHEDcJRwFQpU
yDzEPxG+6Ew7GxTpnONj2U44IhGwPdMxmDLQ6IfALOQr12G5SiKwBvL0Xf1lQ0HwQJd8UyuQYLxJ
lcPQMRSIuBrXc5WaHTSI7Vzx913XwubHGM0p9kKqdRQhZZrvbzLtC0+1Ly5Ni/CKhwRT9Z73crRR
mFWjcjVuzNOXlCr6hanvmq6MYynDJs9muvqpBTT/MadIoSJi1RVqy+jhiwW5bHf2AcIEezNLMg3e
8hdX9C8FqrYdTMO9H9peEkrLniOcsoXUG8MLS1z7ghikItyP7XvRT4m5BAeX+OgL+G+5yWc7WUsk
GB2hxRn/N6v9kMSnH0HnY+wZGwpyBTcTT1pk7LuEPTJSp/dGhwb0iN7FJYFxelONn1Qpvmv29BrR
U2LRsHOozSrD83VHu+M3aYQj4A85RZwyQJaZsdg2+J468seSHW63SOEyxdcyRgle8781eeurvBed
jIaovqBYan7TlGL5FHoX0ycPcm3S4tnzWKI8kLwrX0u1kZt+J3GBsENeK+VXXzWCSFcjiO3Nn/lN
MrbD2m/RlnjYzY57SY3ViZEWmZwcYdiYLVLY84ZP9ZB7kVBJwLYZQ90g7Il3kD9Zjx7flb1jhfE2
GBACTJlc/l8EI4XT96q7SRK2jppOMgVonBkiR9zdbe6zZlv8X4YYx0Qj07tAQN+QDJnPP44AFDQS
hY0FZfX32L0ejahSDkPnQjMltJ4cVNGaDKOzfFPS/jN/p2bj0xr6iAYPoGOYBB/43dGsN1ABYUlu
DJ21JLmvlY9pSFoOaOFIu2OgvlG9JBTKIbCq4R2+Q+y0jWJGP1VXhbtbWYvfG64WfHyu4acorgkS
OYYJj/1aMqbBs9dIlyPMW+Vc7oCIAQskqLEiSPLXrq0olAPJY7XwhjTEcLIxtnc5d6Piis6+noYW
QBY7/KYGxWbv8u3KMZxs7DaW2UE9GZCE/cYHUNVGTNJTA9nQ+F3rqkr6JI3T2LpzBSqVyMGZ+An7
qEZ0b9bOFDTCM7id2xGBjPldzKGCFGEr1hKxi6d21B88W/0EYHxIuaC8Yy6GaaVdaNRa1WwW8hZV
wtx5Vfu9TFZnQMQBQMeDzs4Pvib+eVFh/P9tEjt3Jnmioqs04UtkHCy6UpU4p0lOACqzOWY6TDqw
ztXseMAbq3bpel47Vhp+xOF1vOw9q2/rsQLo4J1j9lhDoU9Rb67FZ0+DAOz328a5Pg8DcWzL4NQa
ZWs60jvTgON2W3xnxN+enC+m/g9dB+zFNHlly0PxPKlEdpztxgtUyhVneeD7i6fpWrhy2nTprr5J
aMe7/ac1uJZlUGELARnSnf554wanXA2B5HbbO8td5OEDwwDrvS7SO4SucwHFuQplI1mdgt43NUYA
bwyP+xtAjv2mFS6Unko8Mhr3VTzWmVVbzZ843ylHy0OMT1TV7Vvu2PKkFeGcMliAV15pq3EwCun3
A0T3bf4Y6RxUrfDOlvXymjAX6DeWF8nII5I2JSapdpUO5P8zLn9VRfCdFV41wV2orkwkSEgmOJh8
IHVN3iQXiNnMi7j3Yjxcciftdot20/drklNtyN1aL/d3AYNRwsYzpN4q80AMA0YYCcmWYJqxVqBn
mMhEMDBuRBBAmb0S/9/I+SfzOfDH0wrQ2MfxCcfdd0u/qHc7UcxCihNnJu8TtbMgAPJTYwyf5WEk
+rmgeQYgP8hj46wpWO6N0oCB9eXMUnYxc3DLTszOdXx7H7eFaLH6iFKLFSwihAesEFEgu+H5IXmo
jDvlKguOgHbS63IlBso0PK9c/rpyRvPOUgh/9yMgn66vhw2g/3oan6NU8jIyuweXk6QRjs+6ZR4p
cOgPOd1GujT5ck1pnwcqIBF9Tcrl6VTBE/DvxCjt0WP92++KNDd4PT60vop4Jd9vnRSmarkhODXt
0Wvj8X4Y8cg0qU8F6uRYq3qGDx/TmIO42EOeIyhtQXTav2jb/MJp3Z6xpgEa1aGhZRwwzjQjD0k2
+3uSWK1bK7fu8ud2uKUohw3yJtLjbhJwgcUWR/cX6Rw/lu6ns5XbAMY/xS/kVuqTGDQ6MXhDTN+X
JQG0pJwVLyk4DUE6BIS1T1p+oyRncckREmHtYo975eDqKL9qTH6SBnt12SHt3CUhrm7RncDw18m+
OCt9JUH8evC8P4lXraF7iq4PI7naAjWsKqmwQLU9XJH0j6pN3uzyQScGtWTvdh6xb7j3xrAtHIt8
LpajdMoLYYhMW53ZdwzehQXV3rD3to5NzZuwZv9hZYAiuixpKHnS/tLiubiM3eYSoWSAu2dd/Omj
PQXabgr1zbvNzyMvwhwPQcsALIAC2ito9BBgdwURvVCpK5vVMMcCCC60Yc/uKLb++tpo82sNsbGJ
SaRsFLbsC/gEA/5DPOj5DrQpPqd7doGDZBPWoFbhpZ7sclmubo3s45K8HsdNxpHS4lW431DcRrOp
uLDKGMvFo2txtp1kcZcLiAciee3kTUSNDbp9nRrvUhy3ponmhUIA+EhysluB36ahXLMw8wGl3jM1
maONpuymWgIOgFq5q6MKTdDj79Jy+gakWcsIZdjOr96l5ET7Trfao1pOUgF+gxDCgv5axuqyelKV
P3iZa6hKu0iHhrBXKyO0f7MCWGrMe3ZSbL00O54Sd7RluBqx8WYHXK1L0SPVB4uJ5wFRXC0RS8SU
cXoa2f+jqEDyN/8vdjEUPbN/IfYa6bdtJor4O67h1MKQOl94yUw2POWjmsblhsBJp5zL7aB00XSk
67LMawGPf7yiNL5NxGAO8WNa4a+6JkhT4gv4dBsfb1T7VcVp9T0Fat6VIT4PnliPJnLEgvkGH27J
41vyODsq8DMeDFmiHX+JZXoept6LBbQbOL+8tGD3XAD3UfCRf2dWlzIvj1UYddKFQ8wsYVomkcyg
k0vgViO//zi2cg4f4QBqA4hszxDJnrRob3EWb360cgOFcpIH4iXpjIRyxyAzfOA5Srg+iPUkjL+N
yzldXbB9Lv/Kbf3fbtGYkyhz1picFHccbuHT8yQhNH0EETcpVDLvZZsPyWu2ygA3qUkbltwcZ22w
TuwknRcXVShjPtGcrKvrcGtWr0ZqXtyxjtOGTyog+WRqa0KQnLh/ifjVbQj4UdwTzFyRlNeepD21
YBJbcIyJRLbFgZ9LwLr1GoU5b6hy2KAxnlHE3rjguntmOMlXFyjfUfByR9ROTbNiEUd0JVnn+ANi
VZsDeu8lE+7pig/vhYqm+0SMidAhnJmWNei+5wkY5+/BJoWyCLJRXiED4/V22HckaJXSHLm5Hz/E
W4tfMwgLkwQ1TdiSkOwml5pHgcrH2dR50Rh9I2QFigd453zXcdPT89h8uncNYoLw8Glg2xrs+vW5
PIF8dO5J5f/k3EoVKilJY+Epn/Ej74F5ssO5TSjAtWK0PHb1CQh21+l+Y5YAH/y+F9ovtD6Dx/9i
lQkDKtLbOSclzbLQb5lv3CYL7K/90zzjQmge5nEzOphqbRumDcfrRLFAE/eXfGLckdjEpGmorSNr
AHsHzKHuSIAyBFWtBuvXqw3KZNx63l05PWPTyiGjA8wsox69MuHVl/Lk9fWxVlSe11+VoLwQFYLL
58kjS9HpIUe/XRE2saWjTn3Vtfm8AOiHILVIZ496JAsc2WfLOd0v9Htltz9lqPADdErVruByFKZK
hgSUftsdUh27h3ujXS1KoDrS8g5myclfUi8mKmamvBd/LXmSqwkfWvFvVdPBdR72t5bxksHCsR3X
MPMvEWIbNbhlX1YFA4/G60WBN0cYIa76bFXdtc7OyU/+hNNIXQHqDtn0xC9+LZvHV5A22s4TPyWK
OLsNCKGTxolvunxUFa1rIKSMEhHKGC02QHlqzT0viHxRtfdCC1+KfqVLhybTafBdY4eQzpihXtl/
P4jT2/Sd5v5nMByZdtLxcv/PHkR9NzEHK0CWkRictCb8vX1c2I24Igf5gVk5F2/jQq5Sm6yD8xWA
RRRoqa2mNZXzKwQXBxfLTsh1P/JKInLhQDaM3xM38i5OivhZuh69QTm7v9JXODjfnFDZy2gk9pCU
C81gGdv8MdnrJ1Wvg6KKh3NHVr26mqIe0O1kZZ4UaRdoj2sp0Bn5WofECSd8X2LWY5z5PF/BZhBi
rD+0s5tycrNjSHpQBQuZfXjGRvH989aMnej7km2cFNYVflSsqWr8AjFSPTW/fZSByhIBvVY4n9vG
MvyY5WLY54YrDYsquF4PrsiGuYAkZWUhahpLepLP2qmyBUrJ8nY9k08bDxMosZ+Y/pWAeLYwTpYF
31T6wxeFfnV4DiO8c7y5ALqe6GUn9OzTDAuf/c4XDIhuBEh/RGXtklIWYb1r048Bkj7ujHFuGZrV
T73isaQZkG1h039fsqZRHKg54h3qfvgCi2RX6aa3hvuouigjhtL+DrnrB6JfaZqDpxk+ycJGZUN1
ykwjBQUiHZ/8aU3PI19jaF5vMKrEMuP7plpyi+UsTuH3qwTa94vBfjunkDLrphj2ySRmbDDQMG8D
5gDH1z9LU83w+vH7J3pFwXpiYXJM0nyeWEtnfKJhXHYS6OwdqNB6nm0id55acjrpzP+Q8zCgYsF0
dcdBZTxJtpedPJdZ5JGZs0MsVu3jYJmn3Pus8TfN0934hLJWCOjItcxRlDM1SvI/fpV9OAbX6uXc
xE+PXbqP7W/JBfOnwUIhWViMZL95f/fguZmPYd1QZOqL7KeoJYCVvMumne7c+u3QbuMB6lAEfZLV
8qB6QdGUs64AxHqz4bldQsfYGU9xUndU0xtol2EbaYJFrjo66vKEkyYtR073nC3k2P7BO4dejbv4
0cmEvtFenDz0g8XqkMJ+rIN3rsUHsYwK2Cn1/0WVdHeaVEA93tfgvjbMy/Ox+sF73J9Pbg51a7Lj
q/wrtW4QsBIdsJs2tg7stpdIPiMVkgCItMtajuC/QcRIQp8cUU8XRK4fRqs2QQCWokDu+g2lqj/v
xOX1wyoiJop+wkkLtzDgNCGmxXhGmGLRw6GD0MQSHQnNWE73YPN4KHorgibAcEg5H2GIeZDAxmno
wRLMli++3LhdBjeTSy8Fzz19kcRKXSEBHxdsxNKj6CUf85TFLSY2iORsZLf2wnyar9arZg+Rot//
rtAvhrkBcW3QRSm4RUTon/bF7273w0Tm6JoYLSKRk8fFAjQ2/XAYN1YivDPQAfWfOBKg3sIyqdvC
5wSXTROE/7lV5tTGzZ9PhglsWE5tcu/0w58IEtzvwMucYqs3AJYHn/MYfZBuYtyaqe16pWtrqGpA
tVx38BbQxTfGwoNtxJP8DVjdGhXIQkldy/7i92o9SkkuPGPUR5yscFu41luffo7GM1OQiMvPwDGI
9tIQj8yQ2149flRddMIiHQb7p6bvpTJgCrlz0qEaYW8tYeGspD24gKgXDR/M5T+WZ15ocgpYX6N8
nvjaoIymXymVigJEM5byPv2sRcUaQGYF4vS+64nlqKwYD5sEW7PQlNdbA0h5N7lFANfTDNV8WUez
cmBoV9QVLeTXaf+QuxTmmj6abra/FdjcQUoT6RDo6Jh826DWMR6A6S7IXuNT8GXoeqGTjASIMT78
h7DGfujE7+olaxfhC7JCHpdJR3VnJfu7sjJkdogrMHWBfFpuqYgAu4b9/NZNBCCSANHbRnfo4sQ5
BCjl8JhAIGEOPrLJmpOXS4eoFwIyvTFKPRGmZjlxCvaqeB7JE+dDVMuwgv16qppmtlWe5Q6PTU0/
yXBIJh4IIcoOANUCsMXDkS3au1ZnMqUHW3WPJ66gFOnRZtfhn2dY4poD3s08o4i1tBO0EsberUwV
emKkHb7eRfHzchDfOit9CVgdQg9FClZTJKO90iRlgVABxcCYNYQr2r/xRTWmlsXoWXY8XIrLGidV
KCDg4uuECxYf4vDpIpeQPllXW23jmERHeHtgaEnWaU6I/AQYM/9YBt0KsotoxFaVN6IVQrgQ1Tkr
e8Bh5bP0C+fYU6hRvBLpBSk8mkmBRXjOotsdx7bpTWBi/yr4iTlqd43qa9z8d+9FsgabLuMrsvD4
PeEkZD7syPPi0thevBPQlCQbI/8TA8YyBc7jh9c7vZFGtpGinNxUC4iTebg1AC2ePXObS2JyOKne
CNcBZbV2rPWkRJig4D8skfoSW/FGDbETVRsIsyA+I/eudnt1T2bAbbaVm4j7R2X3bM79xDpFIsMx
qv/kzNGbM1EBSQdBd7xX/xPTz0NvUonZpXqhvpflbk0nMF9J+d7QjxpR7eg/LT2v/uH8WtzWIQV3
0C8PAMuTd7NXwor2yf0G5/y80xedY5DWQlTSjA1zokhCwtWUGnv5S4OkQd2EOZr0tyQ22fO+YElY
nM5VOMLke6JSNKOPWdboZvEJProc/PRkTSVqP4806nglRrSMv0CA55YfyWCjoZpqJu49Bs7Y+UAS
zUdQxJlOAX0TFSbwLFhqNf4FBkyYGJea/YdVoyVymmNpyVDjxk4fqO91HjIWRlXobnqnTQC8bAE2
V2osH5fRj9FtXn9bYWxXxf9tqp27UNuMjCSE03X2DNbIWVzb8Vn4Ke0i7djNKl9bivkY59Nh9AAU
T1AnF26xdTi1tbQFNz+WVj7QBgceJ3VmCrceWQjQNPVK1HzAR/uWANtMp8XrA6lodDzfn7Rt0VHV
rMlyBgkUo9FMsqs58+wRRrjoNrw873tdOVd/rBVGwvFY32wZwAtCNe7PTgVLrmHU8WV8bgXYelQp
JsRJeEDw8vvm4qkt2zTELUHF+99AOZIU709pVnJlOjVeD0ZqejNcJ9HF3rNteV4+NKvgNCp7jqcT
4lF4YaYU/E5zF6SQ7zYzxk03ohKrhQVkGZWirGb9BkQmz8PG2iemD2BI6yPKFqq9QyFYkZJ1KGE5
qmVPZQx7Os6nbNBYARVoP6Meo8fmKFflSPQrd/coXvj8/iD9B9WuckQETiGUuB1Z9Fm5QD8kJ/S1
RIIc9cM/+9acQDWc1rO33SHyw+NuEI5DLxcEv2xP75AQR/bHbDXH97e3TnWhjuQ0bqkG7wlpLNfx
+zBLM6cINkCMQiwTVRpmbmPiNCCx/CKN+sKhIpJsgPqouzn+Z4i7OWt4EZtkYhFagdU6gA2u77wv
mW2EwhSKEHfr+Zoy5NiD0XsL7hvRH5iOJ2PTVcEwwb9yLy6bTNJj9Ws2WkLsHFWBtMOCBINYxVG/
FcUqp5Zjf3z9Hc42llwX/ShPrGZMfA3awmVupbc4nyh/XUeuwzxfZD1wzifl7ZpOfF53Z/lzAK2b
iCiORwoqLDVfLC3IKCZjSoewWutMkOSOwOkRUvH3AckVYc6UQnUclMwNAFRJcDtnZyns6gjFWAG9
q9ejo28ri9cRh4NItv7Q9eUscTyr8KNgrhIW4rX0pF0S8FWELwLXxdP/qOavT+YxbICuITbKg+TS
r6zq5eXoeH05iLCcKY4RukOeKm077tDihFs0AAGIZjBK+4nN7zyaEu9HT/GLtfml0VEmjXfz7Rgy
oePHiWZ1wdNoDx0ju1zCW9yiTmnKMgh5eoCGXgRmMSgOMbuKJjXpUg+E/XfZ4vwMCf2Hh/4Z2iaH
yzBAx348/l7KaeM6Egsjh4XaAaM9vl0QaMJ9zx7cc1cjZP2DQoavjZNGqlC6ruSx7PhWwHVoMLtq
IB1cksOWvoFsCJBI5A9oUUwJr1MnVJeuqxqH4+iYfFu0jeUztVEgIxH8rgoMRlI7BEVu09r6HJp4
ZGbh+uZGONjBoAJ7m78GHQYloSFEv+A0N73IItU/lR5UcyFnirALosPCSOitGog8tUH3vGmxqBz7
BPngOBL+AS9JB8eicITISI5zcjnd1CrhDzNLfZboAin+FA1kaG3MzdeqqL/1j03jf1W7D+HwOrfE
tUjoItA9HXow2hnfGy7x5Rzg6Wmro7OLA+J7zOhoZ2CAJPQzxeXxGj1tOvSQaXoEPY089f02UQSF
+QHhFjFL9xIMRqQYBn4baFws4evh1V7o4ue9gu+koAdI1+jx8vQR5108I1IsMnqmfmK896NOIC4t
Q/u15zTszpmlyvXWSf3hTHFmWFH4N1i+hSH3puaNANEq+jPAvi5WAbdXUyDsxINqkonURE98LTwe
hpSPyHNRK7ybEKjBWeTu1az5gfiq2aUTUQLiss3+7JOxxSYtjlsjalqSxhk5j0RPgUwfR0fTA6Jx
dw/7/HNMucAdE18wToV1TIwv38ezhaxqV7L/Fmdq/BRyce1J3S7jr/7yBV8HEngE5qGovY0RrThl
/56qznE4VTNLOmCVISZUNkQCH2B4iwfrNjYtUIbDgPOPXD4nay8DqnrXEb7KP9L5OD+nPU0VxRFv
R+vjb3/YxFBnxDfjmMvB35o5es7LkgCNd6xBiqXXKyUXDMiILj/KxhzX52CGZ6s86tRuCOf9F66V
OUvBqx0cuWP4zUlsy40khFY4ANdI6DbGqsQmKkXGH6u+R9LLvhr+bCWWul+chRnuX+qIfxCyChZV
bDMYYMInrAfeqUPq40qlI9Dd1q04PKqIxxAsK7+0EGiyEazK5+okHp/LVzX8NAL3LgmV4oZUmOx9
9Kwib6JJvpLPzAa23GB9oyMXqWUJNDxAcscTcXeM4TzvFgLl5/zYycW3nuDjKsLXRwjOF9a3CHTL
JMERprCJqp9kLYOvsrcuDhoas3b0ZVdPsN/TJgueGEZmCxv7Fx1Kckr0upkaDLU4oYPAT768JVFS
AZOn0qXFihZX4mbTOd2gOJdaylO0By2oe6SpiLYmehQBiLy5dtzTkj36Jy0JEFQIYJyW2/GPDHUG
qcyYm9yVgUWN4C9iKorIdUl7jjGwyNSZ9D4SeXqGrleSMTXfHk4YPBkFwvDv/lNxzHd716+GLSvL
Mc84Nk29k55Ljzsk5Vl8nnVrOv00OI+zC8OUrhZ7RdF4w3QRZ/eXCUJv6WH8EAhJzUOmZyuSqWks
KYnznoSookM/h3sy4Ly3/+OieMcpRlzhxfH99a5hkgbQH5rYXHEaKGzBP5NUFuOJYRtKhAeNpyTv
ZSyO3OBYk8OePotVJqRMvEYNb857NPTBbyiJDFudD8ea7qrK92YqAg1Pe+4vXx4XfnM4LLdWfvVx
qtfdzq+S7zfLVe9Z4oFsbbPiCQWXNmMSIftN00GZq7TPHI4IwZ8lfkR93V7QmFIokkWS9vWAnEVa
sUuxXLyeveU8j+0qzDECnpZ/b/6mcHZj7ayBK+ChhFg9Y75LVy8c5z4ORgXzf+Oaxy0QjD3bpuHd
8RjhWplv+n46aiB5WSrnF51YNUSsT3NK8j2IQ3PoAUKi/MYPTOWtZqzZmIVxZI0hkivQGnv+SGEA
fj7mmegJWbR6snmc2alhGvQ8dNtGs4ghSDwXDuHqcPzOSAyKIYC3YcZ99yQSJ7TtmPdyQiaAD5ED
mglSqXbTPVBSER1vQ7n/F4M5q2ZVu4ldX1EOAQLJF+cUJHNGDPU1GsZtXJMVDwjoh+xjC9HtX1MT
vJ3uss+cQS2lU6hADbcepRwM8dXaTvUXnIYLMx28xcOo18CNcJ2fh4+l+/Wn6n2MwKSZKhpH5/hp
rqrqKnhukUm9XyCsE+ncI6ZEUakF4VvSKwHLkDpV+3OwFvmqR/ZQIXRxU86BUpLffhvx0A7PxN+L
bMPnIHqp5nNskh5YFBfGP/x3W27e3u1BIcmwmzINOVjx7+TjsEuKROJS1c24Uf06Tque5KcDKgxl
mmGq+Uw5dZu3ShSVMmnEtvgc023EXy8BfGRCRp8rdk4SWAuIVjwfIn+ErEETdsAOaCizrpq5tw3+
B5ChUNeYkvEgvMrhZ9nrKO0Ss1hyfKqkZq07OvR6w3WBCnGQoVvl4k9GPfocafReUU0RYqmQ98Ws
aYp0AxBxuwJ6sCuDtEtMG8ODEmwtZXokQUWwtUYrWqllJANE/rk9QAmlf3SymQ/rmv9rSnZBn46U
lyBqGSyWg1GKnY6XS4MbB0F+2jz7Za/rYkY5KjrSzg96LCMpn0MUfZ+WJz+oofBDD7NT4fkIh8aT
usNgftv/ND/IVOuCz6Eit77DR+ofCG7sq/FBj1aKb5XsDZWV7f3fUMs5sRSi2V4XGDR73Mk8CNi6
Q9cpQa2NCsjQfg5uESVR7dBstN8sR1bDMzR5BldI4doKGU0Jo0g1PbqNI0sZXslG4yjxsVizcO5f
7EckRZqauZNTBo4D35RQCmDIyXC8OQs0hxYXs0QW3QNGlhUCTip5LIHOq1KMfQtg4TGfRCFn11QR
2mcOto6vtEJtBARz4MjNY7HxjbWP9TUpHjO6nZzmDgYxVIu0R22ECKqFF9CcKyy3ssqYPLPpnfgM
IisKzVma13c8EldIjHCuBpFRff8zqcFeNdfVlp0MOsE3h841IX4ao/SQLUBDhMVjk+EQuHYnJ0YT
J6CFbHPULZpfvqv7Jv4FoqSdp2yU63rD6tPIofS6sTlBpbbSVaz/vnZ3F8Pm1NO3tFR74NUF+3iw
21FAjXlyu4/UkxUmBy5xll9Mq/DGMDswTmU2kpcx7knLfvkA9WBI6bEc2ShotS98+HYBrYfcUAUr
RjXsalLEZQvg3jd5SIll+lqRjQP6UcLqcIEbAmfqAU7+5UWrU0L31bGix7PWDa21oprrFV4GUa05
WIVpWdgzktwxfXy+91J+5FOst+kEjPISbP2TV/h2VyZko8wXSZhTBJYszZIwqfFBTsFXQZYLgXWv
Ouxrkzt7Xpu/fBz0QO+tamdRi8GSXqihwHL5Rsyn2W2VPdzmGNMWH0HIZ4ecxXcvcfsTuv9mWD1O
8rK5wpImi1MAYOu/ZBC9fiWoPTcy1vbZOB5EWGSUHRAG30R1BhYpNBZHZ080MKUg3hupXuqc1RQk
mYp3KV6UtWjZukdwaBuUEo8QIp2Z3ebnX4TI9GbRBP8qh2SbykGua46PbAakmt2RSFtVAWe6oo7h
eb/RqlZ0Uq2m/9zbEp/iwvZF4Rjvp9zfo8KodIytgh4/XES8l2bBtKwIncLpw2F2vF+zDxKpxwpb
dFK1b5dmvs+tcljJZj1G3euUGFixyFLYxraswn4kWPBz1o08HDf6TgxD+MGnUHzX/sAtwkYuWaiD
kp1K/NcNvXao8FQCgWSfPb1pPHt/b9TMxr8S51Qwo0Ffrp/20xQWnym7SHu2MtVB6dv2Wv52Usqp
Grj/sLPcg/jmSYHEViHlmnhUBDXcQbtSWo26O6ZcEZ9bR6kccXrEqSknF2wqJYtJpEfDKGXvcAg1
Q/fswJl8qqsh08dqbuEH9fCk8vYbOEjHAysekNtIi/6Ra47j9tZ5dfHLy3kNPH1Z9NWIbCxfmQfq
djyfuC+DBlivd6Fn9je7NjOc2IPrAx9AjLoY/kHkZS27GdF8Gle53TsOSp6jTGbZGEbFeKxM6G7T
5Nja1otg1BjSH03zQV2yh+DsgMFo2psSSvGZMrmfM9QaxEn+XCUL74Ad2EB3D4YG36bUGmEw1B7j
VuuzWIaaCMzBSyZX99Jg1ru9lWzWZv0uSCFyBnx8qd6VVm1a+I+hSExjGqpv5I3yGPCKC4+OfyKE
8gcTqJxVcXJC/t2tIIPqIf9pI5/y3qC6gWdI6QaSPsLEq9jY5LI/F1xP/zDJgJ6vcx9bPmheMgDv
Jk1y8oaN/vQZy0v2PKDcWk+YZfNLng66o7EYd9VlyOm8O/izF9K6h1ZqkdUxqrGisDJOx9xad4YR
CYVQElyMF6oW3QIev5paoWhzSHiTK1r3H71sz/P+JTVjvfE1Pzgl1SAxkhONf5rmhiHxtjBNXfSe
BzeLHtqWoDw25ZAXJZW++2S3SfmxXK3KcNtxD5RXd1kL8k/w6R5xKNdlvq1sWEAeC9BKi2YXqZyl
yhTVlirjhk2JzMB5D+ZDgTegs9NWLe72MhffMI0ECbU1ScQH7679LRO+PRiVMYO5JRxnmbaS3hr5
pAF1vAKB0ZsIpbF0Cbez2a05W6I1if2gkbO+BXsB0+TZaFyLlwqQqHHG+zNK32/DzxMY7XMQrP2r
UDguK2TgONvLLIqHaX6318pmtHeWL0mlFHL1jgvs7KuFApJjLiU8j1htUpJrnqqwbbBAAUrXFPjD
Jn7YFpWwInGULMR1CIDSxG4yMMiSrwdBTXrbs11Pytcn16G4deadcmdx1XHJi6J6FgwGm3rY1dq/
Vz8sqs3N5Ckqpu7Ky/zchyjZCHzx810fSqLgROC6iKNBPXQ5vmLMfNqPrfgc7khUfIMuowGc+jMf
ajP+Hc9nHeyHpwsUEcVJSGmH8CM4CAhK7P1rhPicgDJTLIigfVuaTsTAF+wl6/mPGJ4oHHfnoCFX
TzqgSxs8ioLkiijV631cf5Uppiy69+XLu33WMaKtBy855D7RkZbrA0tpHXwbnwqQziPRDMS4HV2I
mOfwAPRwnRMLetychz1W4lfe9Ly+mLwgl38Aegil7YqPivLmmPfl+vTGvonhMTESc0tSpoEhTToc
flpRYiSueYF1WKQIfgBBPcvP+exf9ZgL/+NAF5Km4NSlW9U41sKJSCtWDBS1WE+fQ7rt23nCh1Hf
ejmOchVv4UkSq1lEcCNP3Pi8iP+4TWCE50Koz10CqlyKW9tS2SDst2mnw2XFqkZmT5/Hy0kNX6BU
8FCaKX+chEWc89hKUwShpifsDFBT/xt3A65gk2YZf5pg09Ne5neF5f+/NyOkJKgNDRRAr32BVrh3
lLlb2BWytkpHScNwR+ugtgjJnnwdJfpq/Abx9komGP/L8YNI/VXWip9EaVeBeUkBgik6QSA/YQfj
TObP4k6ahg3AaAISogqVMQ6X5DkYu7SquG/OUb9I9qEi0fuVn/MSdVwJRt5kE6qwRPUoY4bpu+eW
ASqYOXtESc54asPaam0jp4MEkTASP2xo4pS2I52+3eZVIqFdVLOJu8IavHmOsqJVVVxtcc7rZZI5
4VU//pw4S/G7Hs8QhqxANvynhBmyg2h4EVmizi9QYXty3juNB1KtxgXtRs8Knw0yQc2PSbBz6Ru4
u4rL/GHbcDTntZFiHvrUoLlFPkRcVztrgrKAWjsQVmANzSQnlF9QZv9UoRvaslobgBT/mOYkcn1F
CfRwP/wUeZL0L3P6D7lzmpUByE9ibgXqsTQtnV/KaXThyQcXT+vKL+/+EZQuKtOOgay2EpAk9Euo
FeNrbI2CNbRwzL0uaK0vSv5bKvLtLWDx0UDQIKdzVVDaOaIkQLrmB5JqlVRNuIcMwGHpzqxj+7IG
0JtUPYKRn6PoXoYdmjrPl2g/wJNrA/fVpRFn3/vs25qfauVpY2L/gb/zEUBgF05Lp5mf3b3D7loQ
juT5WQ//ShIxwIjhaXAPG7CXTX+0YtEAtniT5JoEdJISw5rQ9ov4KYnugJHJ9+xL1dqKmoSZwsYo
YDUZeUVLTGyKQcT3Bp7gJHaljt9sPrkAVbS9eS5t5wczT3hEeJErtWK6MLWDRt5lZHJ9ktku9GVL
v0XnCpOnXwlkjWKpKOXyLorPcqFA5eeIMQHZIp9rjLYg4ByZqnLzO+BR8XEcZEglt8HGDYtAvVRp
QF7DLjzZsgowq3slgBQB5IUPbY/a0JvfFsWYZICTRBCP0wHAMYvK/yfxrJTFM7/lz1McfeusXQFm
SVAktoJb50n6m8bXibfilEwj8jBwP7b+Uuoh1N2kavY30RbzEv8YF0pEt3DAbFyF/F/kREFLK8fB
Wj9vp4+APwlSq5MUlRfRZe9HRXj0ZntE3fDQftMsWLwo8sbHQSpL/NZ/z/QzHMi+jXlxkltmKQGZ
69XE+FLevZ4QafNA4La01tej5XP8SOc6C8vNq3Wy2H1ejOoL626iTUmjxm41btD0U3hS0pS9+DEl
bmBl6Zcf78AEbugL1bNHUHBIXYax3sjmAD0ysSPcbiGSc2zY4SyMmtMScxWGAdXIEoEc7KQfWkxV
314lhGRISL/cElywiH39pDj3XGW1V85psZTQPWy2iKuHPLbMWQ3BFZmu37VfiFbm4HsuL8vPQvjI
1uCPZzbzrWeXRZwdBfrV17NnLYCtDL/u6VmE71deORKtReYIfVt763umOheu3igOryZ0KyXAcUdE
tMCg+OZug5QrmNqkyneLtDq/q4kIlicSJoBBGumZdVfGK/NuV3s4S/9wTMD73rrc54bdEBYAXc1F
dgvmvbqUCZd1+0ZiOeKvHHYZaX8frrsLjDb4cBApGikV7LQpG54s0YT9Q+PIyEkIKvTtFkUQucrh
bSSAuaGu40URMNMLGFaFwJWUt2kHB929bqP0jMh3J/LjLTVGN6J5b7hwWJ5KrcmUnjw58QVngAEM
YII9m0zUV+uzEvCAZEc/jiAfqIPUN/4lIZ+2gI7z4JJy6fIRYq3lFGN7tlYqPJSB8eM51fA0cMOY
bjBQMSMnPPONjrrjuGulMnSKJnDZh57DUr/3dbqVLzGEoZ6nLbnrCcSR0wGxSnmv3K1RgRxrQfh9
DbfGFHF92PiFFZPzeym7+CuhQ61H9vcki6L3Vt/nZVmiKuzssL6fniJOKtLp+8qBbby5JZtd7yAG
D6RBvhMD4RqKLpHOrSrHRQgnrTnL7uzanxFWKrzKDqoWl0nuB2jnVH93NEDzSyIz0ZV6MoOgMN4w
eQqJv5lbp7lTKE76kW1GDOiFVzzHxUYzeM3VqfKU/IqW0njPkBpv+KyAdySy0tKvy4guEsUUsXDf
4buiwmamu3To13VpIpjv8DDQ7RY1dxh+kvXuTdR374hfUPEHrLx3Z5OrY6V2VtGJ5qqSHacXG1sD
ltkPg2g5EgPo7uTt6VFc7xVmoZkUhnh6nFs3V+x+kRr8UpCkLj4cRaQ59zWrE/8r9lnOYAtwYf6V
jDU8a8bFqO9gTrDKnM7Y25yoDmrOzu1P2yn/Skdb653UP7uWP0q6BIeZvOf25kvz2yVoqb7g5PyU
XKKkxnui6ieWkbyaw7c80D/NDoor9fN/F7GFlQw1FkRvy+TscP17CH2CEPTD1I5RBONof8vvoTj7
LryrKqw/Mcl29RYXDkqApDqioXQgyh+dwICtekzZPepcMhyB52a6nZLDUYtXCmMhNl1juHpMyhxP
O5NcSMznngHz0OLHJeHdr+3sNDUh/weCKvnfzN/AWuFgKDoMHkyyx2Kinq1mxiQ1FI9bFSnYDIak
P8Yx+xBnKGW27ELkEZPnjGLDI/tnmEvzACvJ3mJ7Wwk8SZ7/1u89wGnRNLkmVNv1Z6p8ROjT5ftJ
JvMoYFLIN839yTiYdCazRoOz7SaBGJMfUbhIuKYuYxpCrJ7LXfWKW8ZMRdnI+4u1UiLccryueKK1
z3BRZ9X+KGz60Twl1ATrzR7qiuhsg1MXjAmqscbQKUdXY7a2fZj4Mto7kbVpyn5Litxii5CWfj3f
1HIjHaHMshjG2BTCNLV9QmUgMtTnXbVnDd0rdEO87c3x73zfDjQzFIkU0l446FR1MFflxSeOv5X1
LzvjIGtcgYdITY9y7HL/n3TSAaqlgyYf/EqcHxOdCeovBHQjxTfSP54998NEyEvkn432AHxN4lCP
Q+mjBsNyEJ522knCw3tJBJE1du8G0OmTruoRwQyrWtmyuRfbpYwvSNEKtCWzXYKKl4bdIb30zJNr
uGidrwpWJyS5KPJGz7707qhAHQSnQdu39uS6aBjRXKHFqH8CAQ0ElgnPhCsNMEc1Gj2OsJnbSRQv
zQPthkxUxxsq/kOA+TAnpbKdH0c5QDI0XbtqjG1aCSi2L5TViEsb67rR73r0Cc2kN1jTJ1+aMRAY
a0SD4Hi2UwqxM6KiaPu8Do35Lqh7ftjZTt/Ehu/tDZQAlgUYGACe1uv/A4eSM7g6iA7I3uWTIJfa
9Yv4UwtWowtQ4VvVkEmDySdsLhDrF2srG/qiV0bA7FastNBR32TD6EjD8Xq35MRGUm3cmrK+SZq8
h5R5F4HZ4QNOJSk/VEZpma3u0cyyD3iGI0iwIrw011sccah+VIIHDmNmPcGf7x15E3syakH+9Wxq
wT30iqBpgjme6GQykJhl+4jF9Ag2bESuOwtN5Myw6qQXYkEoEa5J9bsYYuZIgzxAjfX9yy0Xfhjx
3Zqjhm2nDj/pYnJSf4aeBXQin5j3wuIxo0icP+ehM606zKnO9lSCEAvVcDKOk66D+s05bJHKR0Nj
3ysBMqJ+hA9RGYfFLA1Kl50l99OHPntYf0SAk/14+cjjyx8vJT3zXVidn9vkYmxQ8D+fZS/6gDet
kgnHWPu6wP3PKPfx9RCk8W+2AQ09pcI0JM1WkN1jCE60FmiXjTrUZuHV9lbili2VVwoyi8xvkiNZ
m9rBeeYA2NcClUkT3twKjdo9HMRD8ksF89zhQsNLzBm0McY+8dxRbmuOjSPcbWzsQOsAtDCvSrJt
RHshjOMxMTvhnGZ9CDP4AakDPRFTX9oUuYPgAOb0zlaBL0QlhnPq12oPw+P8RaYSLYg4KNBSgh8t
6NElp7riBSTXorsAubgUtvluLG/laXLicdpJ5h8dGeH+TwZwKPCqioencuogyH7UpO0xE6wcrjcv
lZTXKKJE+9sJ3jCrziEjLHR8nDzAzpYSMEuXNf1uyeP9YbohIbi/ixlBias5Y1U7r6gRwi8LfFVF
JYiTX4o9uv74GBxdWHnI/FWMWqnSW3rwyvraeyrNkkKEcSOLMgx8Cu4BpfEhR2peDNOw+j8Rc0/k
aghbS7iOqn4ekYz1j2y9UwxUDdSGqqOCqP4QsA/FWiVOWYeeqOehuPD3yskuJmGHe+O1iVMNrVrh
iS3zBXJTA37jNFMkJIZ9atJtGjzZHszGLAAjYNFz1QFyrD91Ato4ZSl61eIr4jGp0CCtRoCjp6ai
1lefLbN8Zh26lNIj8pK1QIphi/RjHof0SCrM0/QdDCx3LQdq3m6M2bTgxFevHWj/+w09diaBEpEc
tK9r/ER06/7YRLKKwu6chIeevH8oj/slF7nV4iv5A48lp8hPikQ3MkBtDkpf78aG4xwovoW5Qg+K
7xNtHAi9Sp78BPiWZ9HrEAdRa3lsIdrLfwrFib/q65XFqPXfA8KgIbHwOwDO61416PistgxjulZF
MCnC5G2QPlupp/0a7uNis8yWmAaBerozU5FWinqIqkqQoru722KSZz51gaIK26tT6ySyfvNi+NJi
+vnhCXknZ40xU/p0EkxVK/gjt/2WEgck0O8a8fen+erSe/mOyHBLWeDhsCPyieKjrrDBzFziTxj1
J4bXaYjYfkHfHiFwfkXG2PZG6oHA5ruwYPrK4oEj/CbeC9U53flwWOFon8EjNsrN+IuB7jGLw35X
vXwO81ryAP3ngFED7EBzEIJHe+caEhFlHVIfipce78Ph6pKzWsaT/4/+a0tIkaGMHCS/THQWymdX
sSQVfLCvcu0ZrDZTi904TCFnfy04uNxVNP2KA4kbmes8zMsIZEFKng0Wtmy3JlW/P8MX5V9GsQNQ
06Cbuxffa5YSPe1kN0DaXi7spO+iYknvK+AyDdwt+GOFL+7Y9IQXmi9/sz/eF4T9tv70lRaRgsS7
ecDKb1qq5JkCOZMx+LN4fiAjVSvswOoQSQ/aIR/2+lKWtDnC27UF90wjh2rB+VuBJf8ipbKbJ8OD
LgxPBMSSlS9y6ub0kMbBNhXK8ty01aGTRK1mBbVBvZWCTy6AnuiEBf24/cM7yUgkBo8d72e0i+nd
PbPzt3OLCNz7HddVrJecPdDGtpXzVJUFhmSGrCFZJb3huu1z9jDAHDDVANb1v3APhnRwU/0uc0g2
IIrDGiDaEO0VV/Ak5Vqe3yt+GQafkVmBom1McPsdcdnjj/N+q3fjaf92RvE7AHK26f0+KuIWQtxC
E04L2OW5Im8b2MNo63z5xg8PJfha1+AbLsW4AvtSe5LqlEdxBLpLVdpEmufq9+qmzj52HnhTwdZA
f3dI607ijmvsLwqbIW3Gy6C/dsz7WxmxgTLg1/KVR2RjwnsxX2CVvgkFicdYHZbq/DUR2LlD/Wot
N1n3abJ549yxyXt135xgRtIDRF643Tc3nPI7JlovapbzH7g1ia2Lw/h338hvWf+m4SB7RyzPX0bT
GYMSBYvk7el8ZYlbSiU7a5YVgdYGUR2hPW7nEGln8nY99iVDHfciFDskBPp6/UmVfc7z55T9oqQ1
JDrxcULYQzO5puElZk6OEOCjP1Bj3eAp/am9IJ6bbX7Z3cHGAL2RohBoqjykogZ3wL8Q+745shfL
3fG0/JYNOlocBai7e8sMpKpWPuMxj2t1mEypkrzhsa+TsJSk2WiXq9u0pHzEXCp0Oo2jMxKfHNZ7
YwzYsWDutbJhIKgur2OcTZcfNUl0GR100YDcwUSKD0mCuJ6is8YBeNjNnTK4nXngE6MFaobKnqP5
bz2MLqXfUnuyP+1qisxdvjsVt5ceZ8gfwehzbfvR0aj+uUQTG+5cZJtDs+fW7STi9uSPsckoHzfq
sDbM6OTIITlre76Wmmz2VTaAnUKIdHGaMdAssv1m4EFx286rfi01/vTQh0s6agSGG5uF1PaNznMs
bjAOTKZLf4kfDdonrL355V+1KgxL72bD2zDLbisPNZBsSl0B4F6S1bkT3YwomzHV0sI+zCkHqCnL
oOyTTdGeaRund5AeRefNYDYgAVKRgHRJ4fPKm/xJ/Mop0zFUw+lgctwQ/RyptY3Yu1a1W1TmM7mB
ZbziFWBKZnpDYIarjzjRQ5nW9O+ZjedgC0V7tHWJ+8IpKToTm2C3kjk1KgFiHqmJRez3UwIUGK53
0CVdAZr6LfI/02/0O6fjN7tOaIQsOKiGgtCymcD7yWMMctgmDxlQ/99pe52S8EQfNsXrpMt6g4OM
Xk6iNFuWs5x4aQblWNwoUzhCzZc+WAIWw+E6P/NWubfVqQRY74V2cupbkrfvpFOEb/SL0QaGYIoD
YywrpNJlXTUhhyWlolTlykXlv0eBo3pwvFPJ9dIbnRtpK3+IrCfOw7142EzYkHakuS90u02TvByl
r2prZO8Zsf01gbwb9/D1/Ilz+u3Nk7cZnEe38s6PtITcmll9ajFkxSM1KmYpx9Hck5QwEyLa8rJc
/w+N5GxFY7KSvOnBNZRcNTOLDwMa5zxOY1TZ9efD4+QjKoAIF3/GmxLBxFQ3ae6h+DQxXzV4+U2m
EELFbtyUHAymC6WHRsjcdm3i6Z5jPTpWRNzmB9cKN7zRAFbEl2BFaN+V+eAOG1ZZ2RhCkflG57rQ
Y/lz3OeyfZ1fT0KDwLiwKOYy1kU340luElymjjzeLk4LZT92pBbCyg/YedMvv5mes+IwEniv/hEH
PAnWdY5cax7KWdGKpWeZ3NMOltJiuVQbVrm6VdRh2Ln7QbZ7c+G++UsfHThIyh99i+A/SMagtJNN
9Cn/OFuXLeiXiREp5Y3IGkKaEeoNY5Bp1/lRUVAQtvMexHJHgM+ugWz8a0s+ngAxsMz2qynUiDZQ
I9qyxLbi0PXx+eptIQ2b4RIqMFbuN8pIMYbIiliGjTYSLPhzX+6kM9F7JBI00EwOwUnVHmbO7ezD
c+p327pzI7pQtKX8C6Ji1JyyBQHmdsAHGZWHGpAMGUwoKfGUb+474ZW7xQ6v6xcILiGkncIXGwDQ
O+jvWt+W8u0iNUy+ooCHVWgDI8ZNA8YhZJR5XtaQQ0CTOJDZWYXPmwaFz53w26EHRlWDZTTRgVGV
aYcASZYC5cXmDrYao9ym1hoiWHv76I5y1qlkOGbqJ1adLLL9Rc/+ks4uHOWBJqbs2rNp3akjzqt9
fcFQfFFqUQil37LrH4OYXkysrubtU9+f9Pu/p7CCT+EYhVn34hpjw1gYCk5zwz3kliVz4qefHPE4
3Y0ixKVfGgt2HfKWFa0UEIck96mukLQgXVufxsPLnLZNeOse7Yf+uoUYod+o7oyTVtmB0VhFJMnR
8C/dQyATBER6nSNGUjCttVMksiB+A9IfU3Keez2urs49p5pEVZ3oklEZ3nLF+9XlnogjeupOl2Jp
tEISSpteGP4ZYnj5E1fiR1BIAO/MOs3UtA0yeJHOkTUFqAGYrGU9LaVEcV6kyOIC7keWnFW4kZr9
elWDvPXd4rfOixCs7M6T8MXmUpkMiQmHOx3hbxea8r76ar0S7ll4vsYKvgeucHv045aZ/u7wMf6X
m2eiidaZxU3lgm90/eNK6hpDkhAAQ0D8PZ9E3REGmQeX+PNxYse2IQNbQlfulM8CNMVUH1N/mqSU
RklihPpBeBTjT6wH6cAHsmPvfvO+v8pw0XGQ5UqkPu+7Ht3Y8h7DuPLoOvTHrr9Pm5rE4rYd7qNP
D/5MQyZbjFuIamnaNdDT9f0oJigqqgMmBkc4x+fjYRgQjZgCn9rzXtWpA3ut2U3kava0hrDco+jn
RfNTmqHp5oEfv6jjq3NcJt5eNgo8Tdi3IO0DJ/5EvZbdz4zBKY0YzKE1+ScXDUKAYH0AFvjRKzqL
lik8zFM1XAZMgZotMHfzB2TRE+MFafSKgI8qKtbSfu59xBFD+EfcxQ56PaBRB+K2bKtoptlHx2iT
SFvH2AgL5SuZO0zJqVnTY3BpBst7gPFS56hnF8qIW6UP60fBBql56xY56fRHqPNpFdDyzX66A4dW
vkpDaja8fBGHrGSy/mLe2dZftiMavK+tQ5083HqNYX/ZbENeW1xVuUgP6S+VgD8d23KJGAeqciF9
pOd9umatdqkOwisOzu3E+Y/u8ymqejsCUCHezuj8dGhlKo10CSboMwLiaeCM3AjYS7DDN7e5t3W0
TDGA1vek558BpZd3wQzZ/H3kyv2t96Qwm/AqP6uAMYJcnIq/e41vsJz+lEMsosgQJIOk27yITr9Y
28j2/FxSNm1xJNZYQs8ooTPLAkoewf7uOxjl1rnzyUX5Ufvmp8EENP/MXKsZm1IoU3gWaQ2WLWdL
uX6ICV1/vg38r4xSer0X/AVNHmej9kKK/ZhD2SiLOiN98Zf61mWywlAnYOk5MVm/EbEuYwTYrfqP
YdEqt2aCkmmGeluVVViHQH84C7AuMwegxIUwP9brfiFalQgVYePBBaoXY+C7fyblv1iihbx0//fs
NxP9oPdRxEd5y4YlxSKHPm/aFPHo8VsFoyv0buDHkU2NrCryHSYNbo93pedPQ6lTaBZ04qydKwo9
WqyYxaHRZSFTSDmfhjoJWpX1Zu4I4MIwpwBO10rJKj521/2BkR4H9hSpBmvBhx4iNvRgsB0sJTfm
CuSKEc2+/7EY1URUG6MkHuRntlmn7Xyo0Lg4KZjrGhTtmjnSqfM6Mn5KaqnIRpKW/q0B1XzGV+4Z
K71QZzAvfbzC5/R/jSQt4nD9CYscLb1dhKNHPWxHvE/2qH/xFNlsidzkeYXRPs0CzNZ+lsFPdJqM
8m6KkvJyhb/3WC6fhSZx5vBBQTU+G1xWrUMyCrneTaDSeSS8MSZMvMf4HOCifAAknQLDIWbxQrwS
QtvhADzouIGoMJqpZM7qaDpfe20kDVtsgcJgS68L0NC+J412qEZ3+QrgLvLucLohKMjCLEzHeTxx
qlmAHfISnSXBdkIln6AjJ4OuFWYXWliV7T542S200Xz27sdfH+wXDM/nabLBdpmFH4aA2SdgpT86
rRV1Vruo7iPeVFkQUab9poIAabIVJHZTtRDQSxvXO3R4/KoDFSOU7reL02zSO6YgC4bz8D8TP2Iu
vi2EbVmdeJguXKw1WACYVCDe71IEgb7YDn9t6cQqTNOxlxx2/Cfgl1nR3iu2zRyJbjZyY9C2KdOj
Ui46rDyPwotspIPLR0wpX24EYhJDjnuhT7uxRM0LB+VHi6T/fqCsWC91YZnukYhcRm+cuHPCmhAc
iuxm9oSXgEOjhYuanG+gw1oC9MtDCLDfY0C0RUdX+l9/KzxsAtycfjWjMMToaN0Mga4r5azhOGC+
D5QEXBa77YFfnm73ahcWJo/LkYqmcoWjkR3L67v4DjmgmvkVgF2qSSEciAm1YhVGpnwmA14U7D2C
7hD6XtME/iNlsd4ns0wQA24dmGjhhE4CH6RTn5tHqJV1bD9bvjdxtxW6lTdaKTFf+oFb3LGRKfcZ
ZiibO+b3JWB9coLo1ZhaDK5m069+UbtypLAOnJbRkDt5MR/ZHTtxSTSjfqBSGcTB6HplQsl4aC/A
4eE1N2czWoiDHtib7LotG8kz/ammesqIiIrTgVkZ1OtzqlORaAg3dfT+FIwyqdVIXShbJyVaTRtF
1n/kALc0NADpReMptXGPvFL3xqsDL4vU3N+eZhrHXCil4eRl4vlm9adLf34EuZAuTkyS2YO+Sglv
uL1WRdNjj/TfLSr3swb6fxjGTb/F2NlTZEThEgznGYj4NtJCQ74qci3WWaH4aL+mKsRIbn0S+aHD
oVPjFbwixrPoL3A4Oms+Qeh7cBT6Ry+yg3b3GHj06RKpqOZGeWYpHuQngsW38bcMd+pK6AV0hyiP
uUI+BEef99dJjvz137UTOrx9uQ7Bw195ckdTWeWIcmzn0Aulyx5mkw+lEgjK7LlyYd3XbVrVdllo
uHew3oLoZDp6qT6AvIwx+snVS+fsgwngcYdsymfyx5cJbZ4F71+TQmzLCPEmPvoWb3ek+8FsCf6x
WkUB6vmNx0f0PjjEuabME+IaD6GPbMDMGEwuidp24G5lW9TsihufIcv9WGwsnJhQBwQscQWzDke8
2t3Z16ahP/lBoVKqrrHQqncFz99Rzdb1CDq6za012A98PEHCMa9Pfg362ixbTiXB1MPg3wPMTKbH
K0thhmnCGEf/a+BRZWC+O2gq1ayYb+15m01dqv8i9UZ3HP9yaC5cXKAj6A1aMA5Q0OrKnfRbHQ77
BRq/HGWaz5qqgfJyF2RLx8tcrWqe4LsHXRPTSryt3Khkiw2VaGJa22y3VL/U4OebR+BHY+FhmFbQ
Gbm2Rl2kV1K/x3AREwChB6d8sDAYpWk2Cs/adQw6O1DfHi/J5qZ+TnCu4Yd47MmTRkNNdVrqLTwx
iu8CQ2zojh69QAwu12/gR65F1Kqda6qBaG1Wqtzw+S1Le8qKwpD3vTgD6zh+AqnxkdM4Se+0A0Ow
DDnSS2IFTtdrPJuSHNV8wXbeKzMhwdjDozjXynmgWY9I5gytO58LfugzwXYNynIBmfX7l1mpxgQG
Yu2FSnjxNgF6NwNSE7HdGfxNhakDQ18dqM8x4TX2TCliqkXXWX2z4WzJrZcCP6jeIetrnunLX+6d
2Prs5m+tWPEH41h+KWNtaBwTozeVIG1UJmgBxoWdUv9WNCsy406x7Xw/Cz5pYjdEwjE/nNRltCCs
aew+6cC95OIuu9EB+EJuAGHtQbU3+M0sFE9OBo7BBlY7lKDCJGVsckkWDx0w7KQVdGRFEhXKcF8u
LEYNgpDVMMUs1kuwUyRLjBJIB29cGtR00MUxr8MJtR5jgNnRU2NKOiLDjogpfiSfUCPCx2VkDdTf
n03UntpMZm2orZ1M+bND3h+Ym9rAai/PGWNfyY2vSpFKmJ1bOXcUfjQqNoJM8cM9ZS+XOpTzGT/O
E2R3P3wsKPXRkkGoP1BoFQEL3ezRWZVs/HWQ3zh8XipfdxffuoyDC5ObZsC18YGlS8EfNil3+Ko9
CJrgAqFd5ugS/YqrVFLgFQyWflHrNThKVPbd+VQZl5RpP7v4xGInWDYbM38NHN6f5p4vlfM8Pnk8
10xiPSw5D3BAymQho6bEraR1wY/lQLcwVpfiHZHBxUx1PIvthnnRTbHpMl7v4/D6qjjz+ZNNr06f
JGjK0Dqgf7/dQxmtNhXOVFFhtopjXT9KCu/jsEb+Jn/amFKeRUgNFtFtYdAIMhb3pzXjdo8Abi5g
pciM/p5usPo/SsCxNzjUKr3xbpumh28oQ+PoLNOw7BShriRmnYDGMfk3ddgKOoqTI1wvFT14W7TW
cSttp8eoupi/qXnvDtyM2XPnHMiYAHU9SP3b0V2NREBwiOGkYhO84SegVgAHHeSo1hHPAXp+7DSh
iFnMhl85AMw1tfELPkXd/rpx+wj7LfWXmWXGiaNUqavlF6pVqsDRpNHN+eZNUwhqwiqytslZtuJ1
WRmDseybzlWzEuwmsCHqVioRan4wCX4saxYPr3qiJ71NqrhiTi5Lm2exIVMwjQs0v+MJck1zOZyU
5o+CyxKgy7sm1VRuKX1GeeyQC/oQilXQSXLVueJ3sIgzsJKdK5xkjrkwtJqPA6/MkDFjdIPz58O5
nWv4XWY7vga3krej+bGl4jlt9LOqjjNmy7bSmkSvS/gHv7OgeJPGkXv6ygT2ahK+/A4ZtyxGCJIJ
+znlMNGlvAd2tLdGn4Mm0PIAjS1GS1fVecxkVGA7fwZIwNy2z9iyzkaYhBSNtzI8Zp9gC+1PW0zG
wQ23MdHdIag+tktKWUdMlDI3vLmesM0fyt3rggkxW/IJP6W15RQd5aFCqEsmyZ98tTYneMnnam3o
ijtJGcIsn99flCTB3zLzBON0aSpOC/mR8ukQf+IG7GY/yjdFjfTC6UJ1ebR3DxV1wg2v2a8SrGAi
A7sDcauyDt0Q0OdQYmf5lZhj6ohEVszRjuakH9pzmiwm4h853VjInzG++lz8wQfPo5bHbHZG9rX4
FFxN4td40VK2rnsVM8oerjMsMUSi/TAR1HC2kkh5Z9fxbONCt8BmXDjoacwYKaYjjy/ivCgjEpxd
j0hZGTsb/ILUmFMy9gmOICj1Pdod4qy/7l1i3UYFV7m2BhpmtwYYIb4PmsJr61Mb3amIQKgn9CDV
S6BCs0vzqyXw0kdI6twyPMJtI8we4e9oP6e7Pu3E2hwgwKuB0S3g8bmR+pZlzwE09OfHhnBelc3h
klZ/rBvo1Utjk/zeifev35h8YkCSETYjBWQWsgCWv3J90rWkiWMLd2eD9KZGPLLU7fTEVLjU+0qj
JnE4r3tHqFOPbcI9ZOHexQJO6yRxQg+WDIYEq5FTLgGrXEd3AYKiuNvPxUaB5DYtLwzv/10zVbGN
ub/LybX8JYXzyNOHrCuxdB1vp0eH/cezN18zZRdswKkXp1Z2CxTPODk8kQiGrDmtBxvBD7Lnmrwf
OvVQZW0YLvH5VUqJ5CNODDAiI5/aArAI1e9zsRQPfhzuxLsc/mkSS6+nc//SXtyUV1z2GW/5zl2N
siwt2nZW5O54cJcEUzsuo7VIuk4of3NnjPHosM1k76iPwh/IgNDRP8NwL9NHYGkeXPDmJHHsR6Zq
45Jhxq6jPB/RrlHxBHHaZXGihw52BqCzhKCWM3eqPjSfSr4ADT5Rlb3oQKU9ThKUUq3Nf7k3sICb
IZb2bdV2x4LUqOD2ZUCqwpjLhNNQtRFpW9mkI2ypQuo6RjzJKSztJxMSWj2SBLxBZ6wp8VR7JfWn
2SEOM/69pZyxcwLpfMfiD12Dq8W8xhd2iUAncL2x/QWzENF7VnXOmvAZVP0ndQED+1pUReZ8kvQw
XMHJ163wVcn/ArLjov9TrhY49CnCfu2r4LmMmblvD7w5Wyc3YxoEyS/s8jX15Pmrwq1x0dmHKBCh
SLrq/EusYcVvx/FycmNxCZ2cJh93GYDsktiGn+iTzvxBaPn8VMYuKqLpaHmi4qYc/INoX3KHuMim
SNAG40juRVwAT8rvxXsodJCGneMQPApWngsxWm7s4lo1pMUKhqNJ84mKB0cHubgZWHOCyLwkY8C5
dzcWltJvAni1Pj7JpboYgHyCCRxgKELIHcNw44iSAXZw8lP2OwrrkDNtQkm6YbB0SQE+F1Lw9Zmq
C09FMvAEOUr4oWjH4wRIgKSBr06M114HL/CmG+pOOQ3RKxbnjmjxV/K/QuOHXU+AhbjTpzFZnl0g
6Yr3Xv4l+rAKf992v0NMEc9oO58QTDR3EPbW43Q1ql/h09zdLB2RkYjXNER43VXUV7qrpmyLR0Z3
ECWmJgp8wQLiit4UgGNzpUOE1mAKmOM444Vj4eo/DpuMGYtCVOwbtECOiu8AvtuOKRb0S0Fq6+sG
ineBj5e0hq+gyAOUApju6RvXoKWQWA4O8z71f81HuTpREeW+VNvDfV4xC9Kbk/mkib95djNDg2/v
EhyFRhgfOz/9JDR+kcZ1cNyjWErgVNtKZAr3H+KsaeUTueb6mBZmxyl4x5h8fIeKM25Ognf0W984
djjwbFrUTzGLrrC74uUCwpkIwbNEv1YaEOsQ8JjN+67prt3esvIocHovqVSXUiVSnZNUpfkXOMn7
CS5OILvd/6gb357p+GrzqfTrkBFnYChknJBCKMQFxKVr5nnNf3bIc4kZgLFJVrFJp+A+CKpW5EUU
PlOpxBEVqpCDTk3BxljXt2bbw7KkL1pLabh3OARS8LzgttNXKjf/6qmki3MPyIsU2wWnrLENC6wr
ljqVHpTl2FNyyb8fFag6Wj4Nlx3n0bUcuqxeCEitdtrxMfaiDiebYZnE2oFLgOnV7OdusS1SZLmY
tXj+NXcevb7F+f2LuUZSmrxmDN5Un8W7QIYUlPHcZEqjOLFyLzxJ7mP28/MEGg46T4f0ndicEVVd
8S5BOKQkNG/AVbdrhJ38C0xEEb47WivTxBxb1bCrv+M694OKRhAPrOZW4SQM3MMt+Kpy44cZi8yn
8Et6mGaZfu4gAT3/X5ZR2nFW5BXJMx7e1PwNQmiQst/TlHwO8/N3yjQDER2imLyONO72BgZE3OMV
FSHofj73skxKPR92oUEFIdwhDUKgJFGPChQn7BuH0BE6oETX5jPe58dORX2kDLi/86zdkR30vMix
m6ESE+2wWYJ3QpsBsoXlcFOWooSLaHD53rIabw5GZuDPrSn5qEjzKpdmNNMcPWyga84DWj/i2ThS
fkKTXCV3oims+3F7whJHlnf/BRhLmDfGvDWO1jUsV2gj/XTKnZz1fiEvtJ52sVcL1aZiV+Wf2OLI
vHZzIgTSOw1VMkDPRnengW/RAw44axRHxgOGjdeSgbu/+YwKXiscjcJUV6JLCzUj5SooXCO1ky3K
q5bw/71JQm7cnfQInOs6Q1f7B7zc3kjau9OGLfi8J90rwAIh1MrlKnKd7Ze15JboTcfjq4E2EWo7
mKyEu1IeW6vV+QEeAMv4kJuYQtsVn9d+IFrHFIBhPCIpVlwGL7O8KrPnb/SAU3OpOCMRuAyR4ILp
mnFE4SEhitMKJaB0JFPVl8mKvUXZfZxVT1X4P1Xqvv9+HzQHIWr5kmfiqbvyE6swCHz+xamXipVx
GscblGUYqxVBeL1hSOXanvwqe5RiUqP503qCgSYxsvjw/YhxqBJU0jIWH9DG2ab50Iynb/7iDDMg
XPV7uNxtqPFE2Zz5SZaMbGEXCe0y3wAKkJ7UihYXg+UT197tgZSWkthafwl0J5WzrlTZg+kTEg61
s9xcAZ+LDIcziAPaWJQMXiDC5b5AJ33Z52c4ttJTQGQBamuWh1kc85EVMNwAiZLV8alrrUbP2m0L
oq+Ag3MNzbMCcawUxXk1E8Dnd7f7aeeKMPtX+u88Ao/43+jJUiCw/csXWno8wT9SBJasccwpGvER
euF84SRTOaf5nELFbmPYxAy8FxLXQNqTG/lmBupD93Mij/kuFMNSSpfrx4p7Ye0Ad0pG4vSaecCo
9f3ZBbOcZn6pWcxOnD0TZnDEFceXunbRuvjB/hzBzVqyQgPphfKKYN1dKaKWL9NWV/vuRHQ77JAM
twb7khoOUkHMddue2gmEFvyfrASXXsCYGTwFeH/eCmrVhhtsUrybMMXoUJG9z1tUCuBRH3P72hDg
CUadVnrCWQ3o2Ho4x+k6V0jMCJI63/ZV0P593ZL+5ScvZlI0WOobp/+Yhqj9+O2nZOVPURNYSIJc
ySCu84uy3QpmOF3Mc7G72wJEvJtQW1tnd6SQoNaxmlxlMqkZ3yu9fO9h00uZKCZxxOnYRDauOe8C
5x4orE9YKZcJ1eREHDQVqkpID4uuiw9RWwzE7XySK8op/CjDwgIrEqGzv4gc3UAbToI/4+YPGx5I
VmmHqYbgQtur5t81BCH61YXpt4MdO6bf48RldWNXRVilyFSGQVhXIj+ZJzWK1pD/9EaxaHD8qQuJ
xDJpOdnRLI6xmKjobKV1NLYpYfznf2zILctMAoZZYo+9LhXzmtYPBGCPsEwkWpxC/S0PT8UvpjyW
j53fPyXVKfc6cKlRIdYPEB+8aRZjDUVSkKez7ZQcuxXTUrsW/k3+YGes+CFhtfJH492KTXquAR04
peW0P2fIri0aclamzcDiHfTeMnkK78gTyORkOvcX3ZFelvCISwIsUGMy/TbWnskBhaDcmyt8xl60
SB/zTY33xekYQo6skvSQM8EPpRKw22brzpIeXohNiHxDEptBsvOd+a7d5UWngnzr/CvypbGQ699U
98WKRgNyYTEnRkVEEHOV92KeKZ35yXeU+MStXgJLO43pGH9qVWBhCBrRuw786zgTOL7gSBkjdf11
kYUu6NWT1JVLjyy368C7VCKI9gIJdfzYeCkoEei9k4vN7e+3YzKuv0eI+/28OFtIuuQem2cjYVre
L8gc2BY0KAwTn95SKYs+pcKslRBDrNzdJAH9yt7Pmlrot4I20nHnxADytdOt41e1uHaTL0Np4EbM
WTA59rpd6mGDfEloPjGzHdh2I0vdzoUQ8Ng/B7tNO1MP4HDM/TAlkuidH6oucZnwJPMEghvYX1pB
7+HR7DNaQXwEqrQaRrETiL/NkNBHmEvSsaEYhBE0O3hTfWeODSmYAVX/+l+bDYN/sAJEBG5eho2h
YOAJscNgn+ZwDzTp4e+gi5KG3JkP7l8LJZBKZLKHiNjX5iJxeaKDqmcl0Ufm0KKZPAz4TmBmDTa+
3p5AgTkGX7lhHmlP7ZGy40FMZfU/tpnR0flp8lD+d6B6QWvQXgt0M875/RIKJ5QHLdv+ro4p9MNC
ZNZjzqXA6/QZtkrvl8vVt5hyKrmYwKg945gduTqqXGNwRwKYtuREvVaN6W3rYW4QDbdfSu7/FOTP
N183DnokQ58VwEK9oLIkJh6cCPVuOrVRdul3cbvsn/gfI4D3uiM1eZSo9ltc56KBLRVwY+iQwmR4
uIi4zqZFlqpqkhd7GYCLIOwVihBbGC0Nw2mYZT1KIMOdtTetZDhHdB6b8E2qm8ZhbWkYE+dOCRlt
Iddj2hKEOEeES/aFbLi4JviA8i9PHsMgKKK8G/rNZ01J8jqbKyqn7rjJOVoLXW7HYF0eJZ/G082g
5FSDLocq/H3htaNffO+uwykr2pCK6RE9dtZX4g/ilvVjzq3kQDZhrudu70t2G5NY3gLyAB5JTFhS
x1rp5He7uzhNrY8ZrKarBOTpThgLEe7S10yVydPZ+C8ikmotsOxPAvfPV8FIsgWZ+cj/OHXI9GRG
CaMH20wsFwXFH2b+6mCjrJwQOB5nb8xlS5/OlH77rCnzLKThhJKmB5I+B5Ewj6aHVtGn4EBPCVzM
Ash8GoQ7wVVfZSAtL/J9pC6rkYj/u8gKfS6rPNmo2UiP3s6uMyzcl9Gjv/ddS3OAFQ8NsTzGQkPB
t7l5WedvP59hSqCPxzuysWVrgebyr6v7nBwNjnt1gk3pwaK2ChAocODYunIWLf2kAhViklxX8yrh
P7ecoBFOO0AZ374LJIF5JXkxFRGNtm4Pk+yVNytYq5D14eFIlNQ8hNGX2bo8+rVD49ZboTS3rZeb
bj/36odx7NC8O7ys9qgDyup7/27jrzl6Hi2j8ePGZKlQew/RTRj4kUkrUT8+P27eWWchDmNX4u8u
j2Rq/F+yCapp8YZeF9BQBdhXzRqJfftAc7No32VKIbLxhYcpaA4ZCN4Fg1hS/MbOSHRr5WLRmSMd
RGrZulIVDjwuW8uJmcrgky0t7lSjvTuzRF+GGFY/U6VmwVAsAKS7hIPE/cDv/Uct7jrpjSSUL47K
qX8Ne3Bppk3qFBDiLzLmOSU5LerfwYIviaBs29HPExX4/bf04wjVnjcAcbhoUbF+4/TRuh1GYwO2
/hrREyOssoKqmwLq8aL4GrGxdc2HrKuMcr0Dsz/hFdJH+ECkvMRXoX0HIiOgumNtKxHqPgLB7yyc
s811S8lgyagZ42zfDxkjAt0yfLtLs0mbFbbsuV1oV2duBJwBu6RwPKNZfp0g5PDR50ADF8+jHKTM
z1yiqE/QG3XE33TBBSaya3jdQ92u0pvcevP4gXjIr7gQcMgGuZUZ9orJZ1fK4X/ValE667SQR7fh
XJcqJzWEAph9earBw3DtD1RlYmyxr/hMYmrukmHyKMNovoGRpltrbz5KLJfmgUK2ZpyTIx6jpvNV
TcGj7iNlbkfAj+Rc+r9RtIqAq0XT4J+nKztrDgQE4vozPTxMcWAQY+8XZRSLU1sAlU2wrUOs/gwa
MH07KLF/Sz5qdxiXZzC7EIlMhG/zjBKpwlyK/0BqNXpuHbhptC/CjbXw6t0bZXpShIT0iHwdXLn2
jsTqmvfZuMLVSw5fbIveoDZFV5wk7q+zHFu1GKqkIvQqUT4JFj0CuVbOo9ODWkvVG2iCVb77Dzcl
lBbnpfDv3mRLMa1YpPuog2FO3F/hGymYdD2Kt1zLTEA3FXyWWA8A+M5BW5AZa+9v8pkWpvgMfG/y
xvDlbhrG2IiSdSz7AjA9zFSObGlwJQ3b3bwx9aCBjcmDaFizUo7W2djdtr1LbFkdmHBb5XTQcSwq
SwjpDn2Kq0woGBk9pODg3+2OyzF62wD9stS5mMYioDcQIMOaVHIdz7atXo4mSDli7nfrYJV5S+Gh
9sEPi+meOvODtkQimSVnyKhG4oxVL8MImQEo9lSDWAS8hU6gmYHVLwafSZmbfn/u+PzZsb1ioUqz
BN5WuN1+Ho/N/LFxFemMv6spSwKyEVxH5OzFC2QYkefQm5VYwxuNxCv0TxvTeZzlqDn2E2Z3viJQ
Gsg3/qyxF0UoTLZeNi4bOKf+lO7TyH11wj3k1+GcRpagpupkpeaf+Y7whiQwjy7SP9ZUuWu4l//g
b4vXNvbXOwykRSr9f3FGCGccM15ZvkkKAMcZ8ZGoAmR6P14ODcdX/SgdQVIaIXGJjlkMWr4S6Wy/
F3WBrXFGae/kyJWNJuyHz8MKz0csiuofDk5cnFhYMwR83FdIhkhQkgFmm/yvxBEynLvwt2BSpYzu
4DKTjV2Uk7HXleV3PPtzYt9pYPqrQtJZYwwjkmBvF4Te2lRHbDB5fbRuuHvFFAvTqL3V0Zitouf4
ez1LRQzkKhVDZOxjrBJr3Or+zCVqiL8lJJ+lDycFgtzFngokAFSpaLbWys1nrlwk5BILXyr8YUWZ
LZQDIfZjTGlLv6Yv96vrPKL5cyWxN7BkT1Ts867/WLRXIYdXciukqW8/KczDEkfRXhuQ8eNUSL14
fDugQXpef1RK5t6oYQ3/3ggXy5wp5DhIZrYKqDPILZqaOkmfS0KJZ7aqa16Y15C4SRJFyCJjyZgz
lve73FpaMPMmHwOcYWnCqaTskYWHfLi/IkwbyBFb3X7ZNCYpU44+hzcIyAt/sAtqC7Wi4eQFsbCj
z3YMjFOli4s+LQ+Ae8aSGo9yrnwTEJw3DhlKi72RdVWyHMcOPRPTPwmxicg1k8tDDM4Y86eFrDu/
kOLaYMKwI8iJWNFVrntD1RUYsp397lzZd9dBCwb/etSRmsh7qud4zzx8ge/nHjEwUM41ElbYc2Fg
7nzZMqb3L0IQtCTIpjkH3P3H9r6yyQPJ1GpFeoSq71qPfhvuPKNhpbQKfgvcRFDLEQ31KnXCUw4c
dEFs5UmcSIrhBTOTpkNpXvhUdD7dhUgLklewLBqDDx8t9jvF9acIGAjmhxKC0nUI4FueyocxpLup
mABI23WUgk/7k6wUxK3JnofDs+igyaKgN7GPQlFkRUo/B2Ag0kXN95/5tsywTKpCRnQJtr6HVX2Q
H/Y72vljCSjm+DhYGK/cADp+wljX4Kbwj1z7CKLtbQIA6qfHHmPVdN7vWPM8p7Ma0n5971159hML
O6m4qtxLbDRT2BXVV2nU5/li1l+btQF/8gRkBjQkSqJlQ0DVxf2ur5tVPAOG7vzuYdlWpMXEylhw
mcqN2tPdSS4bcROEmDb5qBtk7SnV+RG6p8cZGDYXr60tV2L/x0wkF2iIC6zO3vIZaplydJIIWtdo
8o19ZdbvP+gjtE1HN2RQpmIQNFwsB/CviZlfaqs8Ckf+YNg0gqOy0OOAHbdC20eTqzWYh2dAVrvw
r58BlCz9P+2EB7hoLkivBTVpQIwYSHgTVyy4o1REc985BuCW1hzpAOgTJaQ6xPWUD3R9zqj0qXxC
EOfVb29l7Cku/K0bEuM7xSV2oIZ4xSedL+lc2matkDPZZzOjM+BlRXdnG7Pfq+6fi99XqfPxYxhD
6KoBf57flwVJWLMeTC1RlzDt00r3fsTzjMFaEI0SA7l/6/pqil3DOYAul5R1WwhJB9f4S3fgmq1l
eHms32m5Wcnaik6T4GpzB4V95pEuZdeSvD6N/4Q0Q8Cv1TCASXcCfBALVN1kpT91o3QNy7n/Lndn
UqBtxg0VbYW1TmLtnO7SF3ZExnfRZVL/7M9tjoPIPYAi+k4bqJElT8Oi9pl/DZ5Tm95gnNZuogQc
EOaxJxlXsOywWnE3ojJiiBSMD8WfsgywgzfZgVr2i0CcqIWnb1SfAFSpUy+YxhBbdrg/Y3+bKHng
bSgHR3yr3NEWk2Fp1dHINTVYTfVzlPsnK9V+8zvnhbDM1aIkMcGS4Au6G8z5pLWusaTxRBXhQVZ2
1LNDZ8KKamM3sAQznA6xixhFUZovbDBfwY4XMlHSdRUL+H5Ssxc726iSQwOp2eKcBaEhgWcjG3Ga
8NwJS093cUTS2ZnDx0X6/hel+WK8LVwxDVc2sKD/d0GqFzPvwP35GE9mDxG2SIWKSGnwjdBH0Qov
MRUq6pPH0A9VHdkW30G3elQJxF722kZ+BJTjsP2axHutmq4OeYVGriYih3grh+VBCZs78TXav5J0
x1jmkrQxRhAbAsu2Nf8XUGfdBtBi5iV5HOhfLjpgOCmoyauwjfvFcFyPBBojZ01E49kW3KJBw1Sk
1JmdCAr2HhqCApao/Fc8fqSOdWcRMyUB3yNvIlRFJbeCZL1DAuShlcYDNvUr45UqcJJs4PrgVd6J
Zwvx72siOTdNbmF4CnGaWQppen3Y2Q1eYCLOG89wNvdq/qZU2sinDiQtITzAshgVieHWfjFGk2W0
HHet6epzsbAR/yM5I1HNTY1hMRYbNBNSjxIbgvnAlvhoUwcydxykrHwNVOuxVPzSU3/klXXDUO6c
/vWgLJYXt2cqKOht0sXyASASxnnithYmOoLNdg+T28a0rmsZ2hRZqnjD9tPjhjWFD3wueqiv3tvg
0fkCCJoEFUbNjfMz3Q1uTY50rQ4xn5uHgTtwwVPOFdxg3bujnWsQk2gKRqSg9JSVbtWXzXQ7Lmdm
52JleFD+inSaKxK4recvBBDq2Tk5BKT/TMq07ylxYqQiVE+vWpMNO9rkaMb6Zlb+QMA+UtnOwssN
rVQ3sUzExTSJ6TLwdExnmGr5urLFWFelwwFwuGoN2tHx7lEL3N/tngUzvdXcupHsFynfYu/vuIiX
3ZkLnKi72sDQbogl6mjLXlGAj00Z9m3RnDdTnTyE9MbHkcAv1ELkM5ftxuI8uf3ews0NFI2pEoh1
LaVMmf3ktjPYU4z+snY8FtTPcEbNvSfd44PFjo0wmaDgSHjGt7ivaEI4lwgsePyfqnlx8u0tj5++
4KfaxQH7wLum4yz+BvJWfVXX/WJbtUStUIjaut53sETtDlMpI14kfsld+ilMX958BQgE6mGsAwgL
sTA8Pq2CpI1FVCKqPfxs2lg+y0oqMVLttug9WDEyPuWKhdMZwlu4UhOwMYGwCDwxouGuMnDfSVjY
Un1D1eLIR7UofqPVYiXS4DUTi3YE/5/P9DWkgcN/k1ZvwmzIirtj9ATvuM76WoL/fqSMIKgz0qO/
5KU8KMoNOxUmsVMA05p0wown9B3/7ZpW95mPgCRXQo0TFDPfJvx+eBRebFDbGe9kiLst4AFQ1w5M
bddE04WlkQrmUt0EvQZSWXH9ig+rQBTQRV3aDbWFH+ABgqTD7IsdotYcANIyoX28d6YdJqOOB/k3
cFCJZpfdw9XIoXwqHnnEiwP1UTD+yth0YvJTKMZYrvA0tN/0Q0CbDXCd5/Yran4NUQvsv9lj7tve
3LO2jQ6s9t9sYNkCXwoc58rwjR1qZunLsjihc28v5Dm8NuT9OM0hdfgxayPp4BGNdE/LKsyeMUwF
xidB5+ZywLydiZn6bNlnd1pnv16JwTcXQqg0rN3glaUv6JV1HkzuHYBOTnaB1ex20p9eqC0t0Gor
S5Dsxkw3SpKpGkupPvdjFAR/2FBybk0E6/1sd1YEuFdr0cp2MAbG0CHVSS/pzqGRFpM3XZ0YC/Qx
RI5TxwnAkAxACXF7M1nHAIy0a0vOgDGTql8LjJgI8eiptWC3OMDw5euuv3Qaqz33ZP7luzpfTbul
8oyZpnymqRBxn+V05vVOgNNu9hL+Zc1FXB9g+FUtYD6sFvKDGkw5eDELx3RCfy9kUeBYY+bKhAh5
96oi7GNz3tDBHcSkU/AEB9Dzjc5lOGhqcnN1gZ3DEVEchHPVZZzZtrcei3ceZ6p+BYWoBL3NScfX
xmBkVU0/Z+T8begVqCs1Y02PwGeEQUt19vFqKd5V0fR0VnexbNv+iPUTtIjh5trass40rz6PYeR4
UIj7hek8OmVnM97QlApqNLahB3Qpt6zLzhB0aegkONtxFdXi+4DGsazwMaG+kvnS6QbaoI/sZDss
o8o8k757n1AeRE4nGxpqCR21bCGTFo/cy5Eh9WVCd+VVROUtcFNncbcaoM9R8LVq4Ch8MbT6rJPb
ESeZu98afLcxyF3b6NC6hyrd7NX5cFdGRYRfc3uwIjs/AccakZgnxPc8h9OvapkeJORPbkv0AVy7
i5bZRII89V2a3m3JCEJZIRM2k8WkEVyDQKBFdI1giB/8Bn8Ycs3cRYam3ZD57gJJ3+oGwLOOFG+h
qS80hcHZRORZE/4wt8STn7m7o/E1FdQKYm96x4WCBGWZe9M6QJcLup8KeyjLv/EPuw5K+nWgGiIf
EpDuQBFurzdbftUvRu1bD/t2cyPIv9g+r7tQGgNy7BaIWPAgf1DfUcy/55XE2NJix9LK5bRWhdfV
zsFD3M+bDEqMlku0SljRzGrXabR2Vbi0rYNV5XbYOsqvPDLho5bMe8s0IPXD2muwzrNmtObGMkpT
M/gh1WnD1b/BytS9JbFqW8wkJdeS9uYEJzKeFr3BMeBYKkEcJJoBhQj7dqjlPlrtpawzUftUxvMS
DRIipjc742RSSJgBnMInuqX1xvzLxFqbGExioNEtJZz8ZIWzDr2srImpKOfTb92GF5WDxmOQMedK
tKhdwOcA43qbBkB5Pcid4MFZ0wpLjcK/zAaKYF/tP/NeTuTWbOfpcwB+Wkhc5eKgIMcy+brbkTIB
zRTgaTPLgEgJhq1jZcZrVKiuXLQEMkrXWkvaeSq//bRoBnTuFIxTzRExrb1sMAAh9qIvA+0Re1iO
Ed2qRv2H2ZfZ0INa+sxMjaJ1pL2RYOns0MKqUZU3lcKdd2bp9usJtU1BZ/z7xO5tjcR/0TK8/45D
IxJ48manOCTqb3f1O7tjMqHvlzRPACvZRcmTJEMJWWcCo/081Rqgj0BCneBbvwyyDuy5aLqsoADf
uC+2uJ3LHLL18KbaBqNaPVR11lmyZ7eIiMAA26JthYDwdB3KWnMXqxr+byCr+qyx1MeUIDfENlW7
prgfN+59R/TfZ9yLZh416Obbaa2XyaM6+G2vQ3rxSq+M83lWYq0xjYZQO+WCTi8AlIxs2Trqu28t
RT2s/6MQu0dtUG0X9KWTkEmwx90DtabVdKGlMpRlbuHe/nizaHggLnjjJXar7Vw44crdsWWztHbK
DgG3mlPdf3NKMMRwjPmCiHRtE/FrkGSH7VbBtrO0mkyY859tT+kM1QaeFe6sGaG5Yrz8bQUh+ZC1
+yzSBpiH/Nh0BgOfRb1M9jf8NSbjsew5sXbg+PVEHO4b4BEoVBqRENKYX88SCDqZA0lttGvpsPP/
LyoxHljfhqmi1pjckoXsfiVAnoSYhYyzcAquedItjz/ByHUiEpAED8qQAzbHgRjfc5P5qQeSmuAU
6VISrKbS2xJgIbNJtOMDFNqBv9DY8kR8MW9WoJGWkMCO4ovfdEHU6Fl+9YvpWndlL5Fc6fsL0JdS
hPswZQdn7Bm7nXiSmiZuLNdnYDecdyiKeiMu65FHsOcMTVWWzBgp9mDcvYpIZOl9JMBE+1djj7En
79LfqWToMAm9F4q7zZFm5ulBGQHRFlbNzyDx0wNiHWH9UkmZBNTkCxnJ6wymQTN5JD5UjQcYCjA7
J0P2Bq0uULZGxuSBaTGYlIBqRbjB8W9f94bSgAs++s4dfpHjB7JV+DsHN7yVQdAnla7zJ0KWEeBd
d3FtSSsB0Ld6JTlUvcbAzOgMblIy7G7gzaVnW6MifKRskEnpGUJhuSa3CfRS0/YrMLRvYY52K2Rl
Td5iDHFXed0H/fL1qkxMbXVhA6ylxoW029vw3RHlnRpkkbEOKheCymow55SujfxTGKaWF4zgpXFa
ph6MOVLjsfMzBsOYzghe9Eix9nU95fGXZr1FQAHJX0RlF7/GN49XynzaQefIYV6QqEXMK0BiVQGG
XxdspzB9o4vBDGw1OI/u5Jq0S3k9KZdRDnafaIOtRIshLcdlnn+UAIMM4jKXcpoVgSSgGkTSixkd
n86O7lqhTtjGQUQKJaW3VOjDn2HEAU/zWl6cdsOh7quyrOufJ4RzGxXz987ZxbCdPG/Rh5HNrZkN
KwsHM7vJTY4mFUMfTCfyNMS2jpRIC85mW84mEu50J8NGFZe69YH770sEijtjsKEIjCFRdD17hLtr
4RUHkkeRjCBX6FDHx9Y7jYxuqEuEanorF9helzbsF2vkGDFmwmnoOp/Dao67T1mRxAY40hj4ZtS3
f7ABbgmXzSkJKuHpxiBFlNeV/PmcYusH/G0hlKeqgaQCxr9dx9V3gHspgdoq5/WTW1CyghL8X+6s
sPVrDxocH084Jvud1tas9gI5ATAQOWiikyYt/H2gNb0NpqeDlrdxO2oTJSsEQUvpELIi18U9y7t+
jhX5Dl1deond/O3j77grd6ftBpuZdMubhRMKIPeG1me/xR2t/UufFksr/+FZpqpgJzc0/BC1H+J3
KLPri+HMJ3hTS/GyB/uN0Nxi1zswnlik0hH7DFHKTBdha9gjm1FaD8wbR5SD27hCJgSscsPPrkc0
VjwEoFl+USb13yw5RVYg24WFw3doUk3L1FQXv68wRMawIr3itzvkh+xWOUC02i2IBnL4zmaZQlcX
4yWQ3D20qX/RnXSCUYacRV+XpjfxqIO6OO7+3ocL4vPtEB2cyKiC8AkfUGVhtvkIb2uL+urDHG5d
UGxTkcUvbMvk1xdiHW3HEaxg1tgzfLjRaKe3eN+1OlirwB7YsKa8bDmX1wEETBkmkmQa4MnjeCpD
c64K2i55JX4hqf7R18fapsImf88LQZbXuuST6Cd5US8UyI4kU1l1/KXcMgA8kFUydw54kduD7IbJ
0cip2H3wKbhd3By4oZQHImIxvZnrwvBgHLXo9YofmX2XBELzE6mWyL/mdi984jhQBNROAY1opB4E
xcPm0qzQydOiU91zN4PugBNbuSXOVVqjk3yEWkcjGO0n9fYehcUwB1C/fLtJPgHk9eIMzlDXNudS
qChFl0rlw8RKf7s7lwBJlKUhA1OHokGpianCQ6HsIA+Gn0tAvABM1feaYTdxQSN/PrKfZk5UA6RV
KvjcmzYUMawGrDmysfZtjx8WfRhnmZkM4byqmOI4lIC0jw+8vXlmbenaV141+Cc34igM0RQyoQkX
a/Iqlq1oIMnBBjwGbg4ekLUxDt17BPqNwp//hEFOqSd4SW51lexTUy81qY4rygQr182U1TG5/E9k
Zr2oLzvUaGZuARuf6eK/mIDa3q/XgiTxH7HPhA2fZvdLSurR3X/4k1CQntAJZV93Kj5dz/FspQ75
+iWlLBxUnY4UmG/oQEOtI8yqVMefls0ov82Cnq/uoOGBva9max6Q+SRu+jGlbbSy5huq48UO8QUL
D9heu/PE2i78BRaMO6xRim2zMjo3YGujLHjODV9S4acjwqaotujVITUsgWFiZCk6ndj9H7kw+gnB
MT8vU+TM2FRgveszGmdCF+kJPk+bPunv2sEUbKQV5cvkAIxJdBOw7PPvzWQ6qLbu5M/sTdNkN7pA
u4uzCORJTI7cAr8RVy9kquOJOvhnY1ffen8T+TIgbHZGB8ZT0g7NC1FIRIXm5LWm000/sBzNhnnh
Ikwd46mqwgTZSwKbUKFKyY1ArDUQ4PB4MkfDTJHkqRLqdMmWX5lGMWaHL1xcCorp2mG4qe5PO0On
8UBlT/pGF8eMaK5FY3u+/vrVDYW9XWB2Y1C4JABXW2TOV8ywzi/lFMQFVR88Q2y/b4p+1cYiQCuk
Of2LZKU0pSvoCilYEspDx3jN7Hqhs33UdfpCm8TEYAqpRKRu+j0nGVpsJM8NM+qd1WRP77gTnmNq
bp4dhKxOCi1cUGwUK73w1zAaTRSOV8ylZ6xKASWhXk3IHuItuztn29EWHgwKz5+O8FW3uR+2jfWv
JKrhfeT2RazGJJlMGqUotJ9p6fQA7aXCNKU2+0aFfWg/kpGjp9W4vS6vBOSA17IUP49MKoKw4tvz
cTObWCZF963UBlg1IywfUhmtAJoGip5WiLwqAcDHWMp79wtYypDdLunezuhXvGUbV+pArKF/xpm6
2zt8DZi1V+gRVzGvmubMC1WfziIEDpPaASyrk0WvBXRAUyDNLvOkXQZ3k3/rAC8an7aUJgG2Hmt9
v8hLY5FzOKDFgWl/KJQil2RhEOA27NVC+Zfl55GzFb2KuyBgSQXYlfREeN77EOzg4Z7lG1LjZ8h7
LDl/R/mNyPqImBeuUFlCteQoZNkJhvcixUHUM94TzCjbNAP3YBj636LZ9jFJgxeUHPnUbonjR3PG
ZURdU7XrndTXuQJz9jUmGC5133TBGiIDk+Z6CrNpCjpNWCYTqMaBe6UUKFFcrKt+ERyTSjCXYqGq
3qEyxxWVmbHe6ugLYgFUK3JHXlxXMB9NCNSsZboQnJubhtsL3SQm0vOxEjObh6mZMcDrwZ0sbBBi
Utm/H/cGayXYgKlYc26rhEQzyFssqi5DTbxEy8AcyrilxSbNfTEUBjuHSCHHPy1ecccjE7O8NfmX
ljamIiP2jOPGIx5rLV+/zXTSpkWFLkul8ZAxPlQd0VDhw3jCX3moJ0qtxW+BxW361C32AfGo7Zm4
2d+zbEdW8JO8RDjg+QWvFtCPH2tiuEwhzr+ZFM4Ruo55N2LZeI2EhXCE4Je5nvm7WmL0VCA729Yy
Et5mAWbii1PY3Zv2YQF50A5mA4A6VvzrKq6gJSyO4bAScjIO66Ouv3x2U4JVVCKph+GjKxupnicz
4DtNOfKJvi+re6F+Pzv6fuIIVZpk/nRl2UDNFOQZZ9PM4QonIqbgE+mhhFJXb6V1AFPCwVsL3p6P
TWr85EofiSA1GsqoEWPPAIcQpOarmbZBjxMUH2HRG4snpSKPXrasfcZQLkYdSut5I6DwhvDfl/KA
3HG8H0fsrREWDJW/YllMC1JylxKklVKZED3TmicNmab2NBVpgBaE8PKQRUK5kYWtLf7oS1EfToJ5
TB3JcSVF3O8MDyklprtfHN+pwmHp1Jp8HqvCFYw2VLAw07Hc9e/y7//LJygb2XGwPSbCHWpKM1I2
8Kenx/ZXYYONEeR+I2imvYchl8tkIcpn8xqGixvdn8vUqmRhibE4mORnZu+5KlZySLz+QLvDR2NB
LYVmUmb+GBWMKlZSovStBK82TS6gtQ1hqXTEWIjBQQHXv32tyR9tkQTYO3eHnDcmwfWBQfhfQfao
o44MGNJR+EV0hwD2SbOf8l8iR/UuCxr9W8+pQ7KROuUNHou8jIoRhKHkGhF8L7eXvQCldbyyvIl5
/57x4+kYM2ixGfi0skZ04AVZtF7NFjr5YJfmKNtAUkQwYaHnd2QjNqmJy/oly1B2TxnKflBPmgf7
OGYATeAmxXoy6MS3iMWlAxxQEK0bzKk9r6L95qnn9Kaz0M5AmeCwvh6/kkDfbhuprS3FuGAKP6l+
XLohZ2KAu9w0bVQwLAV97ocpN6Lws0biHk1VAbK469qsP314G0cj3Ha2dPEHDNpaXgJXnkEsLXQ2
To0PY4V1U4OQAAEGjcoTtdMUQLGCMd3MGeNhyOZTKKT8ngVJZcadotgoJMmrK0JU0hU4XsWvKOxj
eyg//WnE+Sm9SoFPnsu6bpwHUcYWYhQpN+r5x4zlr7F7d9R0+E4aRRsujWK7iXoA/Y3mbclV8L6a
x9rolTt8u7rcMHF3RorP034DHDxPfWsb/WwYLynbURhmx8aHgVDkQVxhV4nnG1Ak3KYsHms0D2NA
67W/0y/A2px17cCc4MriXJX0CvqUlprcBKg6XtSqh4iBvx7+Rj975m163eu8tRf9xdZIOq9Sl7D7
PJ7sAfx9wfxeLQ3zSNqtMwrSWOU/aYjqe0honUXTP0RAh49CdTiI73H6bHUIHNge4OvnqyclV+wn
tZZfKeNtdNxk8gZuaQSys6Jmne64gyhY/KtwCeStKr3vVv6zo3MikcizyuIwbU9ULb5RDda1pKRr
PJabDivnYXu3jOCAz/KYPnnkW8ALK5HJHuDl3jEoN8pFOhqFFnINhAHGJtaNJZ6Lpwn0EEWo3LGo
HXkyqK+JfiMY9tbFzNfmWQd6fGyoya8R6zEAnVrJyaAcdF/5AA4BBO/z/0t2RFmT3sBPwYKEgNjV
IuDc9aHPk6fBlChRY7JL4rmRmuA+zXmZfEgrGMGY4H3+HwC/YxSt55PN6c9y3UQjW5HijXBOYESG
BhoJioEnWnbxOwdtAylwpEOMby5mal6SNhNXnesOY9oTNcfshsMFyeru8NRNIT3p60btzYp46eIh
MyqOnLNdvaOwiMa6YPVvrArmmpieNxDYgpUNJywH6/4+wjPj/RrYnMptzx/5Af2ZkGV+jeYro575
i/Y+orxRQ6D6EZjEQCobxc3zg9SjWQdckCznYq/+UsEIGQMVpajlGRivy7X44iYByUC3o/s4h+hD
VMKRPXeXHvVi/Y1youxx6FzuJaC0IxTbjJ6jCD1QTchbJf1cmhESqsCN37cUz7vgWDukp1cx/Y8k
GyyUCtesbVE/TCqRAPFZ93+JGTl0A+68gbc02mOj0aBiiw/KEVyBvlHw5q0VHIvJgs6w2/fpE1uv
P3SpGPR/qnFtWCxuPoxlOz1BA3SWBbe9lmDHvplt8G2wrKBGD1xiMO+4bOYYvjRfPXYlOiiJWxph
k4W00Cwrtel5WeEimCG9S7MILy0KklRsUP1yhvrUSdLzk4gvBEASD9eB5siKJw9e2xtq18gfo2Ts
uzt7aS/w9mg7yiwnoqUYWB/NDODD1vmW439m96HAg0kFWUpyHM7kYB4XfJ7mOXy1BPALRRfzOfsR
GJZFI+OsxTcrpxHTBsoPVAeP3YZFY2yR6eS+yrP5zdAp2JySwxfG8omdcPhae211WT3yzZprhONR
aLXHH6t3GQ9nTidI1esMJ5PX2vOZV9XnvwjtHlht/toawYJ/XJAky7TlAnho0OvETG4rlLLl/Dxw
QUBIftbf4OjpdZsDKQr+wV9fOswQbTYHSgaJKvtRt5nGY8W46fA8xfhoduL3sic0jz4AY70kD/p/
ZHU06xeUQwfjEzvGk8ysp+x2RSmL2pJYZ/OuMEutzZrYQ4+c6yzj44fPn5S2fo5uFXNpvB/azYIx
1fmr+cnWjIIcewrwH0+ZJGldQNmNico6AvhR6wH617bHlyjgcm86nwR6eEuBoWWzBqecI3V9yUsr
nLYR5Sc8Wf7BHulhNFjKmD/+evW+OcWyivRN36EKae2/BXzgrJIgE17CS785FVPrEDBA6rb2IJUj
bUSTQxqPkEpBDehOog3j8d2Bt/D2xW47DcNrwnqdU8VhLtTNrLsQiw6kK4CT/WudwFWrT71UxkF5
cC3f4EnJ2dzZqfCbKdFYt9q8LmrTk6Q28HxjvU8X2GrWf9a2pbS/doF9+TsrdtYf/sox1kueyZpu
0Bu+okZIlK0QZ5j4sRLHVU5wskyuMM0uAcfseJy44I0EBjZU8GwqBxrEXpBEHjQXYuH2obKwUNQP
xB2Vntop2KBhEuEhUMd69DGjtmO4nhcOGbwgQbVVtXfBrwBigs9znjXzWHviXNnJ0fqffysaida+
Rh15UJ6uLXAIQ1M+Iov8gFsZVNGjK/FGr8dySJF7FwEfXLInIIRPK29QlFV2J+nYTP+iwrd9x7Sp
a6+2X3ZqtjCkvXzhe13Gg8JHwEUmVDsaNeQSu0UuAkE0bKhEbp19yPLjGh4HDI3ACMkI5yn23Zx9
G+PGwCBIv/uz/F38+gwTluvj21TKOkzetKLnIZU2k6SvvMOx+lL5cYk3i5E0OFaWF8/rZKYT1Jzf
+E11Ry3c5w2vemqU16rQ3iUHSzeJAv2X5KbSdvO/o3jNEIHe6r199cCAFnKJyEXI3sTwOH1N/r7O
yW3fd5sTT57ZR8cYMKPz0zD3rBvMHtookqjXpmnin9WBb5ET8ZBYJwqfQJemah2t71COmZvtVUcp
YCYn1jQpmlnSvZtSW+yyvk0uZPsVKFO9yzkLuBC4sKW05yXcdG6LhZXK6hCJEY0UUX+28i2SSrfg
LITvEOgMHPUmviQ5o8lGTGrjjQZ80xPV+JYZWfrJN19wcUZVK+xsmozSI9QUH2ds8PAv/15enyhw
lczXKbWl7ee0fHU3G+Myjh2//NlJWwFqOCgG0tlUNQOytflctcIkCmAhz+BDkbzAeXC6ADK7jBY+
v4Qli5/x/M67zqqX8xD/dRznD27tGpCvB40AxbHiMZuWHbJgPm/cJYwkhXojA+odAJKZvUwAxz/w
kZaEOl3SyrnWWFdVprevMhsMOSBDzxSNphH4+qeuyk851i59rYNaMMWyxpOf7O8KmJNiHHQ1hJPG
fCaFRkIrthxPr4iIba92YOcy3N7q2vo6ycamQaVM5mNfRs7IU7l4RImrVOjC4XLvgszkTl0stNuE
/kSa5juHCKcgIFqQ2j9dA+mrATSmfTgea22m8tiEvuNfNpGaRLeC/fUclne+tADqwGmbStYvY5TN
ZRLll7swNx6XgQ1RequxnvzzI4rjuJR6CzamFcpRtgn1WKDKHCKtY4WNAMWfy0ugYwEDk5r3SUld
4A2LF6L2v2M/6nzKkAoSsA4nrJNyWZhiCNPSYNDP5iwGTqCI+8mnJvUjmDmea7971r0R4ksY5Bc/
nVFFmoKDctqOveCUypojthbJG5Qa4eP4JHylwDRCpVCqDtB1niLF4U4Uw5DjR15sI7m+2YpahDzy
k6vtOMubbWpRNgCjaWSIULLZi93HJl5v9G0JEk69NOJS86Erz8T2L88b+dZvQtDZKeVJvhYE1r/K
mPI+nJ999/azBqtKkq10zvlk5ja3UnzoCyVpYQzFglbcOMMCmAsdopHNUQrwSSzndGUbMhg9dvdE
ahLfftDTqbMZSkq//Q50NJWthOhhBIEdSSI2dLpUcMOQEnJJOzgxg6+mc8AY/yfND3shyC0zLDKa
3NMPPNneY8Bx9oGrIcFr4dvi7cFXhC/o6LaDujfF+Sn+ocNOC/wgQaJy/1qHWIF7kvqaCxh+Ljdy
ct4qIhFFhBMkPS0z6/rEz838ekyR7aBVbfPbOwgiOKGHNSt4x4K+BfI3BotnjcgGU8/ODHkybBll
67Jeu8/8SbvmxsPNV+QmWorf5o6FwDfmb2i016/snx7s5Ivd1w+pbBcbh5h4dD87ovIV3V8KOOcd
mAxo+3qAwwl0ryBzIG4XbOpOt3rSMGm2rxpYAfd2lXYUwEQXtbTDulZ2aj7veMd1ofLtvop551XH
jwx12ORezw1CzhHcZ9ffHkrjy1N/g4jCgE5R7QJSMhsBxu0WbqXxAODpqraiAWhmXPCL1dvTk12g
boybA+3wzJ47cS6GKuYNzEubPXH3PGI23FZ7+ljh04OMLtkJoGe/y8GxcuJ/cI99OQyoAPeP2jDG
7AJwMHSYA5+QTZU26Fto+JYQeHFEAKsMoTupC2Ec6ZjZDrZ7owLHWb3Ihegftyv6VwHyhQSSP2JB
s+nlmntJ/J+M488ZG9vYcxPoZwNBkvqHqbhpXK7c9TAItDZl6IIW/9dXMCwsHO+Akc5LiqoeNPyu
EFUZtc7GanhWMeH7r+L7lR4qlc2Mbtjy6QWkt1R6U6GNczjgCzDwxR/fh7y4XIv8mlLFp7v8Ppq6
AWTC+FsEYID5yu59DTISrwSlF9NRjuN6GCE63koufheBffMwqHgnPxghQxfaeFLib7dUwI0nzKQK
NAl8ZZlBZIZ85MYlqPK7G5O+2D/fycCN6lcdLq9mbDDglM2ufW4yoDRMsSKMpayMr/+IipH7eeQo
skr8+5kdbv6eU4lMVJhAf/znbIqLD+9r8zeXYbTCDw5WvIE15cA/63dBTqF8jLHCUtIA53sp6/09
ZbX/yeLsH0RxR8HUm/jU++DgJNSamGQdsgG4sAQfEecSjiZkXf7+k/q1M3YmwJUUW06DW9vivdhm
9SHMWqzv2BtzBn569yI6VjDfhfR5tbHPntOD+JQiTIg6jqvlrCwqPyCw3mzIEc9Otf3dXdqEtuza
MK4XrAQhcWZib8euEohU7hYG2A4italYrtVjU+0pZjVgEGMyNfZQXbxtuBcRTdIejKo1Ki519up+
E+7qDzPZ6y6Cj8Ta1Ceng7NDgwqBhrCsfwafAsQ0bd1bhpRH2iNg9VA2zzg4sfe/oVOugpRaNNdb
xiK31HkKfM997+92tZI5/a+BcyXmKSKYo5dXLai0DJe7Abz/g/fGNpMPeZQyjkNRFWCKT/5fbcBc
RG6TA/04DCt7TrlgmXwtUpaEpKYltZ89dQMtxMiYI/BFih8e6fw5J6hKU8QH4PBq7Syj/7HiPvcp
l3q3d2nO7wqpB49iiQa8Ts7l8Rz/mBR/fqCuOzN9u5+fD9imVpIoqBgpPLQiA1nMezBo545znrm/
CU/fVdIfT2WTfBFK1uK1M6XiV+7zcpo6TLCgKlcq7mPzWJVex1bvLs8bjAPTtIfg+wWsWMOgOaI8
bUwYnqUgE4YnonP7gfMJ8JwzA0pruun1kkJQCiL+W7lfvBV+rGB+7/QCUEulb6i1KvCiK49snmcJ
SnKtDTEBWJU26wQuv8r4eFcgVM5uw4XbLi4ELjIxKhqPkBWAOmYcOce16T9ciegARBD0swBGWbe3
Y+ix84k6qZtm1dglC8u0e9NIacVQZxf1ZPhniHdElmo519/YD9yqxcniExMlouZeyFoF6XBsmDqP
m82oPhqkm1aqe/zkCfQxSI06psgRWPlSiZ+JvbJFqtBVPiwn0ZFIowtlieWQ7fHF5AXYdlqVHoMy
+3ZAmS5ZR4nz527DdNLK+brW6JZ8fhEYt/iF77WEH9UFIUgS9hoNr8fOU210M5j8wU8xmzgdrvvw
jNFlhgbmDISl4gSwi2Q3Hg6cnCNTuqDupv3pjDzkk2pEKcLLthe/1WqqeFRaPtX00mntXiod6XBK
QJ1Z3bswrd10b2ktCmdHDPGUJVD911lLTQi7lKLOUp6fmRFNd0Vf/64YIbDGPJF8ZZhrIQBOs+I2
XtJmEL9zCMkjtfHc3dUiLUMoUobI6q2Yo42/WoXqlfgFdXgaPCkVb6+nsPuVOSZTfxkaeD/zfuWr
KnYx+yvuo4B1TctsqvXR/x1re1llKRNFmiEVeVVfeGHaYjb4GG9rKfnO3t4HAC3bDDy2wO8EkEL8
J6CW8941Nw8zGnqutB4yxZ6BkUeK2We/F6n+V9G6AxQZ7sTlO3IazPpfNg1XxYIhi9SGKgPNqD5C
rJi5r/D+KaRmiroh/09HWSOQZkXIQ2RqgvF07QVLac2JOMfaMsrPPxoV/jMlUcUkVtSNmP+Nz1aw
H5rv4EBLkVhiZfz4ARoVBPRmOad2UrHRLnla9jF717kwlsRk3HbN+fESFmialDQMsImlBdshMffa
0qndy0qEoIaQFrYX6pnWO9pdHBFc/Bb2I+89IX081fdsZS1Ab70rqUGnV880BnxaV7PSNiM8QTwo
IISofl16WZSPDfG7LcEmGsvsD3NP4gUW88PG/zhop9JaOB+F/FcdUr+dMW/kFwM/6tsbkdTl+tBQ
00ie3GvRyu5BVo4KMXzCDEfTQpcVecXms6IN3lznCLnr0hGx9s1pY6Kxy1aSH6AYb0230xApfGBY
C9kfrr3GEBDXZSRZGVB3pKlRZ4Diw+J0XVsoF4g7cfWMW5NC/JOKog2P6Ga4u/9EFm9fugcmhvxq
mWesyv3Ir//yk/OaEQgjTf9muQmRWtcCktNE0Q0VvDtrRzlxXBys90AyW+BKP4l2uQE/vz4dS9aT
sW/pssHgqsM5XnkCv6uqwIAVdzcujWqDw6JNhlp/6d+qNgtrVBz3uVBarDT0CmOz6iWHGAal5Iwl
udS2VqDjJPzinQWYx1q2yQAKpOKKF70vsOzOkDvVQ9JLevBGg8jUSWNUzgh7xdZIw6+ksv83t9TG
qjS8f7KI1Fb3yXi7iZYtDPVHot85BYlMN0uR5soIdIvbig0uc/FHTfuZn6IdBYbP/ZPA05xXrp7M
Sj37Rwl+bk3sd7d9cAFbW2iLQs+ZkvXssZBgcYfaE4cp5YEhR/1UWjSIw4xRo/dNzPKukM5AhNuN
09DflGBKzCZrpctT6PEJyJpjIqp3aKbEDvsgav1ub8oG0p20OSmggPUGtDtHvUfmWiXcIMGF38Pi
kSVKqxM5K46QLctE0kvQHVo5oupQ8Cc5FQDgXjbSZjCMVZmvZc9o3sQ6vw/xMmb0mqY1KDMAWU58
fV/vvGX70EQ2jGyEh+F7djqO5XvpzipG3SoLB9QMlyeFqZXZwum1hcFZPr67KrgbPbqDx3X6a6Ap
RsxjEWBbjej51Q310K99Vmf6BNlnfKub/ah+GaxBj9W3a8jcM22jl9Nbe80WcD47Y+pQb2hg+CkO
/kFfCor8hP5WxaGttjnAs16D9LntUcZqnnpC3SyPTtUgpkjVPkdS7q9jQHY4hkrcGxRe3peI9GAJ
CbiRRNe7Z3mPXabysEwpTIRvvzpZSaiCk4V5x+mLyVuq7XZGiJTAK8E24hJs0s7wk9cfEzsFtwOk
VK5df8xoGW8xsw7pPkMGXtu4kgQR4f5Tc5teb3DZkb+x8BZkWHBOhzy5qPFq/Q/RcDutkikrS46s
RpbtXQzjMXZ59CdFmBwKXsghezt+fdsxwUDB5MlgGE+WESqfUyla9dIhpE2bv2NJWzv50I30Keha
TZQuBip1HN6SlWCkTTyVWi9J+V2Wxm94/8bO+Qn8cg6tYPaQUuSGTmntMK90DqhTE0aabKwYZX3/
J4Oz0xDigoR/Jq/TYmLHEa45ZRI4ZJsTtFhyMA89O3lKbFbfRlN/5lyIMJpu3iNyYcmXA639MqPF
vW2DbE4ekcflo4sLG1uEd2QH6FGm0nMDR9NYarHxX6ZDxZiUfBIeZreoYvU5hknLnqkMW60L+WLS
FGIIvNf4blw81x7Fjr7XxqFkxkgygXnVPP/4X8iTCKLuX1aisgbet9GaJIxM++1Nhfx+RYvlTgRg
CjaM6bym1wdju2KeMj4OKyamhmoIWpMRfurFYNt7cHppx1sjNCgXARzGJQCYzg2E6mUPyG0DMW0f
0OkmyF0mskxTpN1V2QgFwylRp/teA3XwmDAi22O7UNQJybL3FcYrm0JPwg+9xS1cgiwa15C2vbhR
yVuWvzNCV/ZteLvqOzJbIXpi7xpoCPYgUnHEVhakhrhc5kfTUP7i9q+0xXYIs+KyVLqhzTAlKqEV
4vc682A26ipI/erTw2kf9Q7wbB+CqcEhQSseA7jTiAHGTlplIps48DVEmocJle3aL8zKGgiwQn7T
oh5fCe18e8eBHS3jOOZ7fklw6VZn8BC5BIv5h9sqY7PiVuknZsUShcX31v6jQNinq08sA5MKJRiv
QBsABDcCCtOJWoCsb2ZQa/97OxGpoMhYhVxNjAtyd3ac00lAhbTtZHSQvdsnPbbgfig5h5uro4Q5
y+kpGtcryZKw1aNZrmlBueAP4diguQOyOli7n8Y6KIQWgCqHKGM1uPrDGPGYWEcdlPObV+2ghB3d
TkVaRoZ1dEBb/XA6Pq6q/iJhvMon6VVcgmASlLOvokVm01EVWbkTxkdpN3sES7s0IwshrgmybAF5
HfQPlP9MCl813+lBEAMbUX2jZhYS+bMjuN4TfyapmaI617hGn1YbA4+W5jJtAvuy1UYksf3KEOUY
VzDUO1eXmhSZ/XMnnzJKHWWApwYSGcvtYpLGLKsjtwWoLd8XA3cOCPU6xgtdg7brmQAlqJlRZLiV
XjGyd8CCO3XkSVSH//rBjUvPOs/doLZuuYZYFVvIHQPVhe1XZJ3/QrdOmVaGZ/5n84b6No5iASR0
/hm9cuh/HfRABSZzCNzDa3o/ZJxbS11gsC0CfyAIPMdt5+ROwCpYGMeiOmfMPkyAJZPj8+H/ITxl
e07V2qTML72ltLpDldO/uTSyBG94tBXBy2HHzwd8/+N6Rm8xleM67wfSoqrNntX0FAO1PbbIbqje
Ta9hObGltcHX+ddp5tAl7BPeoH6Kn5ZmETSk04O0yEeNkDg5uBH3MrkXMkmj47gcJuEssoYR2/MI
rbWyL2+dygAmjWCRA7N+R/YJJR4i0RyxaKPxHWFHIQhYP3/QPn4nUjcxAQcjmoddNFcV8bDsnwVC
tBcMcraaJ/ZgQooRGMeI8BWBFRqb9iWb7YoNG9O1o9SYjx3ek7pZRsq7yZic4hBdAkbY+rHg7YjB
Qi5aKZiWiQ5OddiWPcBTsrqKx9BfEfWZn/OMVLaR91mN1mZ9VL7wnVE+aznPj4sPTUz3VT8zlgIV
c66jZQpWpqj5Zu5x5WkTvS3FgvfoS+yomST3fOgH4pLwKH+l8EkFt7F1TDThVw4y5QYT07ECyHWS
U3h4wdzpxo3cJNmtrnJfpE43sOGl6cXz9eqhDFu7dsUApYNHAZvuwhoUB4kXjU+V8x3zEHoC995M
IzMbVWOVWuSsmf3cK6uYvqR2xqMW/H9HZ58jOg82OLv1ILb+WeDWVdPlneLVjA9MyBRddUHpNw8W
VDAoHnjAAOyRFdsOz4SK3dgfSyG38IQ+j9hw3Obaa41Im/eSUU+YaBFgAkdh/pjTAQJgvBaTYAh9
Un6yV8P+pVbH/8Up5d8dcvuu7Jb29tdxA5WjtK5/N85W9YUSkrCL7NAYqL+/mDWPGKMf7n/ZN0yk
Mtl9wlwZ6FhfBh6xgXw5t/A4QcSscrzS0QAf4nFKeFXoyng73kLKp7dndj3KgcF8JqlyPlXIP/Gi
fQKnPl8Avn49G7aDjvxftAuXoBERkEP/IMXHuZ/WaMFIfsEwNzjFs36Hj2/GsINFUsDMPn21yHPT
40uVzndqBeL7xXOx4n2a634aMFegH3PUhNqz62nt1TxxeC7pxDonWQOKG5A6Ioo/LS9nB2dWmfd2
gdPGlOP7V88Tntn7gePeL/hkM3nrDxYhj0/6Oz0vUStVoPIPuKWBR6Z1ZW9cRQk+IWcnUF0O1CXE
6gxIbc/nqsuRNU1LVW52BDtDlPMhMrHbpk9ufqxl1sMZQ/RaMgabdopQVUL4RjJa4pxMiLCOH1hn
zM2VbhhDNu9bcMzZ1/HZb0Y/YipXTOoyiagzliRZVLKWxPsGkqSGx6Uf4pS2s6XNItqgCWoZr/1c
4SWyBNyM4TK/8Isn1JZepUiz5WiQox9wwzkp6p9KtztPSq433KE+jFXEB5xpQ61gvRPCRYamaNgd
VP30x2KYQ8Scf+DTT+Rv3hH/gG6ZsOZtIiW1cUx8yQM7Rzp0CWrusgRFMm0MK7LTviw/XT6TQ6yR
uKxpSpNm6fjtemWym09KKJf6EdVLeB5Mej6gkooo63fRSvNTHCWjQ31cAjZ2qysar1YiPQ50veU+
pa9EGM0+gJMH7zY3KyKUWvilc8DtrGHZl2nQIjwLfndk/DzpKTHVPD5xaQ333bSBNroLaOu3fIGe
z9QIz0arby9xmlWou2JEq0Br9oidw74KB3rGJVLwjxOfZNlrBVKTlKOxypBqqRip3znPcNNElk0c
oFilzVRbrsMoeXmL8tlv3kb7SD/iXm/x7M8qe0Yx/ZxrHusAqBGvlgTKDfnLZhkCppMCocPZOGNG
aOTRImhBPlJEY4F5GYfRba7giMrcHc5QFfaDDwpIFkG+12IzltWrOyUDaZNLXcRFIyRP5HbAjX+i
wvTT4j6xsbMmnrp2qnkw+y6PcRbmcR+P7JEwzfE85hkJAmA5zDgv32BjzGUmocQq1ZNKPZS8n3pr
QPbu/oD+Sooao0dZvLdrbjFdn5NLGubqbBGgrwQuKb0wJIEZjmcUpiJFYmT3AnnDojV3ONBtQQIg
D3DcioCz8b4z2LWZra3rHnthE9myAuLcL403VPgQVfr/oAhaOrd6+yhRqIBBqba7PiddtynUU54w
hDq0UeZn9NsYmJN9gncriuJa6w3wA/txRetgjmaaY/VXaH40J7TB3TG43dJso9xnG7Eqd1wCReh/
9ePIfVsFRHfUj2J/m4OCdpVTHqouv3hshQ0fMiS+0aL7TvAUIODeekvHRJ7Wub2fo5VTRh3+EfjD
Sw349XmChsoR0a1GmwFVQyd61dD0ufnmHZSbMh5fffrfqEUO7jxrvM0lQ8Z7Mu4AHKLoGW85chy2
e0Z+3Z0IpRU/TQ57n5nTPcsg1hleexzOqywVTXe59wpwYq34WcYiClyI2lDQMl+HrvT1hWRUEa/b
VydT1XykqRIek2JvFqFbM8rJ/QA+ioGwZb3UMraA/GSFtOjeuJuKdwXrBfCdBRyJQ2mjtsVeLWTg
mBHfRvzP0j8AGCYW7YPqNVn4/v9e9WeHmupUpnSPERgnmqyXmX00Ef5v3Jmezjlg1AMeuf5Zb+jq
aPTm34YIlSyzeto47NCK+GpUSvnNaG+orQPDc+HpSI+Ed6uJuMChOioD8guXyZD4GXRc9SNUYwLX
73wo/QvQeAuHyDNZ/hDOs5LBWTAn/aGJeU/9NYjeQmPcOz/dltfX5aa4ZHNJdCfI02xDRlC3uMjr
0N1vzF3IOn42b14k8AWy/H1YcqrntbxJjx6l3lJK8YscezUGqixuXpEDrHO+NhNlSmUfRVWO8LUd
oE2vqAu5jKCcAJefi9N2YO1GpablUre7buvxXlx4oXHsNPDF6EalKOe92ENCyZ5/t9OPkG8fFvjB
4XCN8Y7Crark3BhERYnndmwtn79SUEXHUw8dJZsCuuN/6c+WqHXA+hTEQYYI7DA5/r/D7PwRxf5M
wZ2oBE9x+0kt5JmaB6iB2TJ1Ltv/K7hLxqDccIghsGPmQLa8Uzxl+8uEVbi+MzUlU+2UinJFOVoj
YrIVwaN8ctoqGRKQnBp9MuRJex3P9DyD0eMjQhjbBfX7OTWPKpmbktxr7TVw0s00PO1NGZa+FZfK
1G/y42O8ZrxJH6yx6ZvuQvgrjUHPJn+OguLF3T3jpqND74l3EYuEoJq8WGQ0OZovMu85HGIutiyP
uAsHfxSyTfm/J25C+YM7Cee0OzzDZorsAEGvAUQQPeyPPCdxCxH12HUKJn9uE8SUEzac9hOth4of
gxVZGt9YfCjKRT7HrOdqRJNe4gMCSM9WxG34pkx5aCnwJk0oMsXhfayHeYZUNMrg7TtOpp4AEK+y
GylnEV/JxM1nY03aaZpQ9rlBP0UaB3zsOdEzpzlfvkBxECTWwAQFpjcf9wdvkAT4bfo6OOJgmyO8
4quPjqHuJo9DKCyUq6JEhHCbrAFTUVQ7c1qni39jq9lWFfTxx8IyURtUEa7WHxFlpt7N/Pj+hefm
sZUvEHE3kEe2ZK9micb/edEKa0mOKOTXpSkzN2g1ken5jn9G91n6cstU5s7XS6kIksFbRkKzyqMX
a5YjcFmE1D6m5HEMpEbvtYdCNwGCCbTNC7wrdunm7jKn2Egsjv0fdU31nkx4V27ccNtOn0qf+D6S
boRWN5/8fftR27/F51yEruuW0Xg/yGTeRLRsrDeizbh8NrFNDDx7xjJN9GFzgDw40087urEF2NvT
Qy6UYfO9pwe4+qd4ZgxG2Srxyrmp8CRl8+5NCUZSWud7cN+YgW2cZ00VQoopt/5ALe41Hr3Efbw5
lonH0l4TXikU888jut6QKvKjYMn6b/cR2Lu8GWirWSg0aXtC6RXrcORO14u3Udk9lvehAD/uSssp
ykjp+OeXRDJeN3JoRA8DlhLevcduOUXeW0P2asgjdNeErxBUdmsb9h1i1vfb5TxKhABolDIIOxli
gI6lKlq7FifVw4SbRuAh/Kbe8hklrpFEhxrHrcedDzUJb4mWI9otjnjFG3SWccZ+wkzQSde9HD0U
2KdOsUOkat9p9DkYZdODcH4+2hUZ998uo3/3wox+bMEvv0S77sQJz62Fv+b94STIhCq/sCPoxihT
14Y5JgJAehLBkGzGSCpBfJ1DweJpoKlfLB5ge0vrvi51Gx+OE6WWIi1dKxIPHVMb5sF7wFhVXMwz
UCxbniU082TN1PQ5C6SWIbe0z6377ybArV5B0WmpjoST8JmjHJJ5sbI+j5bi1C+iPlcrJv20jXuq
iNAs9LJ7LKndegkgPmRGS7ZrCJZDAz5L22X9PVFQbNG4I51AEp2+cr0nJMaychYvsYBB59yhqSno
HFTKswf+W4V1HBQk4OrykSTVF1zROVWMvsTh0Z3OJpgJPawiLjuwCNnNG3Njm3biGsdnSqY4AkFp
8+a5l3H/XvXPYS3a0OTz+m8Yjx7amJ+BX1aMzliiFZS/QTa2GyyYwB0hdHcLRBGJRZoyWHXBg2Gs
+41kkmY+wtJT+vB872/a+oVFDfMOzqUrEtjCEJX9kTp+G/ds/Q+M2NPHA7ALpLTvJFKrL4PgQnXi
PLC0H8iN3GGjBz2rj+XSJPDkHalHY5VOxpNc6VmUKh+xQmdcwafmG6aamMMr04hR55SAlRIVrgPY
TyZd0lM6iVwg0+N7u8alDHa7hlOWgB+OYfP24XMUcJcdTay4H2iIqUDFTfX+7on2Qby3RZIuWNmC
nPUPoPyNBawC0rvRBITLarm7BkafnLwxjNzBBIWKSwzVCvT8MaW6w/0kuf9arB3QBP21zjSWBdTS
z3f6kOuhyJEGbrQT/JkDKhopce6MH6DPcRHDof5EB6dL1/vS1itWUTejcMrkIJx1dUlSgRZt9z4p
38G1xsFa4gYSQOCGq3vgu1Y2WsRjA+a2XIgNoVzaDZ512FM1HpMFxUPJRDx2KoSUFCfH5lBvX4ms
0Zxo+rJKxryr0JOtcCzmSnKs7YIJv/5wteTYrL/616GcGvi9kkSuT0Wkx+ZntfMzHDYjKXH/OZ23
B+UqFI8ja6tk9jDTXD8PShRIbKDimIvvHRtRhFzMfph5LByuH/Y8fXrG1CL4jRAMr8K8zs+SrB8x
CkYaxNTWUgnpR/RIcMTtaQ2EvqmxHLFrEYu3qB8D5uGmi58Z4MNqaaBNbfjldSM/Jvz/RwnWL0LZ
cYCc8POMjUMzhnWYh/MKQFfbbpJ6sOtpdVaaTJ7Ve7fWoSbIdJeE4SLL7s4hlwzbRUWmb3MvMbbV
Am8cpPS2b5oLA34/I197YdOdB7l4lXnsKeIuYz5zSiH7cf3Ec511gUtebNojTifyrAQI+XNpwlfz
3AVpLt9kMq18W2qiPmZx8zN/D0hGuuQ4W0sQ4ihpRNqzsHXF4WNsrhRd7+RQwstUkJ9wSO+toKGq
cRg3wLfbL5sxPWK7Cb+7B39BFbTijR1q2RieatycPO5PHfUNeAhs32m7ABmHQay2JGxW+i/IKW6W
2PC9ka7Kh01F1B/5MFdQshNK868UWv0zsWA10GqBwrYHfdHgQG+HHmbxt0se75+fytzsMntugl6p
78ztB1ONgmCtGGxbQw9xyESAhj+JkDzbnFapnFoHDXp0zGCz84LledGVWA3vwyYBlsOLfl17IUzk
lAVCE0Gg2/ZmTVWUHNgn0B5p5/EbOrfngkxxlWdtWz1F55kjVGTa+nSfmOm+DQZHcEZhJlkeQZIm
SNnWtJBbFnLwxc3cZMy1ABBGfRz0gnD4n0/UWFPYrh3aUrOeH3opm/awCjcd7Lt9W/wMn0AuOk5Y
BgvQvFfsOsEU+aEocIAnL15PB/tbKqS5cvH9VDXj3f0hAIcuM1yULK6JWF2ODosGP/juqPT7nMj/
8haJsgwZA46LgaqqyXhSNlxAaHabV6WwmhBeAlF9yRgmqRJ6+vaYDn1pI1fmP8jEaTic/H80UQ+q
UQYLvjCqegTa5slTKTEeTfd4Qgs0w4PoLlzeal82skJWfuB7WbzN1toTYbYva5QBoDegdazoBTBv
bIZM+X/bf02jIjVG4wR4n+r1SLCeEN/og9CWe8YJnDNSv4OahtAcEzJgkby+JMRRDfhbIoRuGiWa
spwZLoI8yU2Tx0ZlaQxA4DTzZP73oNtzRRQTuz8iOycv121pCwiP/rAdGcQEN3CzROa8N/I9uSyK
7rLddaRcpxu7MzlPm2jMOBs4zJI+lCkS1bJjXQM51RYhClkhnjdPmMhtsho19mJDR9U2aYwpPm8A
l7lGvdKEcdnNWzjbcugNcxa64vtzhrXh4ttNvforuDVcJcJHgx+NVoRNJXRK8r70wZdMEkqoEZFV
FDpRIiAUWKVP4nAM4kt+RpZlVgD7+o6ajOj/+ysaFm6ybVZUWHzE5LBRu3VUOk8dMEcCWsNrPzj6
xRw4nMWHD7TEj6NIN9j8qSQJo/Xdya8AbW0I3F9d3wkEwnMCilg2P6eeM+NAWSxB9D/lcoIqea/V
mZWh2+pt9YVTnqozQjj/Bsz7kglGBLyUoqgXYwBWFskVWNhSeBepm0/rL8r96YkQarW7M9vapgGQ
C1mhlS0+iQA5DSx/Q4OBqOku+kMTlKbo+2kOTOYDDq5FRi5vhHZ0eFym2PxvuOnM8Nxxb6pPZKIc
7XBAqdY+dJqw1aS6RRgsSe7eu1sYuV6JZpMOMoYTA1WmhGoUbe8g8VVSz/uiGKsTeS3w9oOl9Gdk
NUUofJQuzlrbW9en6WehT8+QpMyCA21EtgGNNMAvPqbqOQU2xZbeIyL9fh9gu8/tnqdIc9ee0q8X
5K7ILEXSaBUBqOuQnKALnYBzioKdw36lzfthYpXcwW/Vw9k2aDS9HHSFrmPmpNL6zmEqs70eyhGR
6htWtuf1xRHYIPxofnXk0XBjwmmG9vqCyXSZAYLs5OgjJlFXyhgbHHeHHYmLxu4gSKFiqLmX/Pmy
b8fU9slLcZe44cK3rHSuj0xZ04+jqojDJROP+zeOALK0Bc7An6VN0gnzaO9NQJGmFDrt97nPLzyJ
Gy3JrCBks9grKnWwiMJ44Wit3kHSF3yWsCHnRsnAc/i05ByK72FVA6keM3REkJx6M9xolxseXQsQ
m+4L/BllWet7LdkvFiB8EN0XdrJH0qmxP9hnWkTvgRgveeevWPOGSA9a1RFXKAET13QfteDeLK0x
5c+zZDc4h1z7zGMtewaeJcAZX+hHUwRy4Uoqy6yU3G+MU55JGWXWP0LEZGJdDQaZgVWx21rDcrzb
jWSJTA+kK/FQnHVTRfrtknvS4NGBXJWOA3bS0KDfM34tN/P1UzkG/n1d2rJ9LBC3lbHQxLwIDpNw
cX/qO41UBbbruKtEpFN8ikj97PNke7h4Ft39bmFa+OUEFubm62ep4858T6wiKW7ujovQxVP4NWEs
JVuNBm03UqXWyITRQ6B1ZwKR15bcVkXhgZBs3yHb7TyLcrUBUrd8QeabY3eQRlsGius4rqYIXmLa
x6IOIrUxNHhpJyB0b5HU6OQQlqP3VLB5GoAbbiVi+WqxoGfIJYBClGhqNuzoW+PO6sL2auttGTOW
cQp1Zc5waz7m13X5oa5O7FvQ0y6kcwuauhJPcAGHz77SPm4baTxdKhTD65H6upxaLP++igXwBGvv
Z/wEoSAj428o51IuuwZJEnCBMhG1eRHNX5RBd0Erp8+n45GnKvBKkn5AE46hBZbq5/VE0jrSUtlR
nhJnoCzgTNWgIZwRBdm2OZTVQxwAKm9D+MK/Ywde3VZnhYiWQRe5vPh2MIOsGH2LNlvehO+UMoHr
bKNbonaORcT71fNbWnftHdJBt4J9/Ccqq88/zdZHA8aCf8FkJpegC09v0KryKDyJIxrErz7fuHT8
Ll6CgoNZtlyjHtmdbN1hOMTMZWSugPvZDjKrFk9QZhPiiHTlhqmzw4p+WUG5HJt1odi7YcSWkYKR
MssWYOdE2QDUScF0yhZVq8tqjPotyUiBzNWmQFfX2vPznE+uMWHR7uNTEkzE4g3MLr1K9DHwL3qI
/+yHnGmJCxrAfgsoIwJhFm6mVdG4yQV28QdYBsfitPT/jUM74qMewmySCDRNhvZIC4Zim5D4Lyxf
j/pS96KQTMPa4SvSPNWmI6RwqE5vlW3EGZrgDHFt79ojhpN/cksIid990p2cSQH4s6JvCO3ePB7m
hH0K1LdYjYwEm66vtULBq7OrbW/RzErb4imzdMvZqpibLsqb9YOr05UH4DGWCVHYfToH9Xk3GSiJ
4fuVAWBVDVrH3WckDN6O5jbUb3YpLDCkOhPSFa0UV+0TyouWnlSpUCcIDVGeof/xjpz74XHJViHA
8NHBIG/nVDUlfC3nZX+DXxYBS0VIE6ZHeRiwppP3KGAGxmUV9UEw45zaIgXAfMSpNHHPEu4BzmLp
EmhTZwQt3lzjfPI1sKIvoswlOMmIaAkpXnKfC4RdXyliCC5fDxt2TmQ80GAOjOR40FB2gWoTXowZ
AUl8YkTwAurTfeFTywm0Cikrs0rLJlj6khGiI/CcWM/xTiW/dw1qkojzIc1MuND4CbhgFi0E3Y9j
YD0nyBB3f/2DqCuaFgmVs8bdW4/QC6tBMgiMDBCo998bpqiU8S9U92xpbSUk8uSAErA8jljXEeo0
0mGUnXdpDX2DlD6R59jj3zlwo0dc9UcVTU8pI6LWon8G4MBfARKE0SAKot613RdO2vTjzYpkox38
s/UWCvFywAILTPGT4G85LxUObdwCG8KCbeVHAkKGHuwu9GKSu5Tr/2Qj+BYW5zqH5ePPcK3Hs4eh
uUPHA/fGypImKK78WQaWzCc2ooTwLQzW1kCkTSJlScnqVCtBcT3vcnnK6eePibWCmKUW10n5WmZH
O9QIrzBV8amOKFwdURa085u/LropH1V2Qk+bt6f3gr0UhyCcUPqGaFudk/QguUKLy2TMPLXKSovV
0mzv+dVbKznyjpR7zOKrCK1WKhd63x68MnQbuQcs17w0JwPv85QvYpZYjpTlEMlKOWsYh1MM/S3x
641WLWC8dMKSr5GwBztlnVM95iQSJo40aiNJ4AISddTY/sgeFTWw9ZnVOZNd8J53yxuSot0nsq13
UaLolJ4Zh9fjZuLgnMSUliCgyBSvrFEjw3DJay5UraOA9f75j9OWjecWvHdLBeClSueMYL8+y5O/
iUNw5RK9iRJ6C6NsafAdy4uid1ZB9+BPcDZA25nEeTYnzH39qYEIs4sx6Rrum35SQbm5alWgiN52
aA6hKWYfWhQLumO/YghFmwk2gaJsOialkpH0LMOtC/D9SnSIEpWDrIocDa3o++XqzwTn6V5912L7
3W/VYDXDv6xpefldSPcBoZPZJGd2Z6h9alxTgHZ4qSy78SkJCv7UK51zs3BKVzyDsWbrC2aGg5TA
S9L7pDrT3d9RsOhg1cBJPXOVrjgbj/Ct0F1EyrwIBF1qfsT9RBs76xh8GM4uq3U5oluRfosBNf2D
eHXqBribjUeO2qpaZAOtg00Bc4olbXCKZuwE9nob/PFMBszCWbnKcuzSwy1FEAvfhM49QeiuMht7
BnjTgA2YBYGmPZfXrHxlrXAdkogxmEwspW+N+3SpibWCrsVzeT2bO3R4HYk9UDb0RNisYiwb+02a
D0LcJ0XCPrS9xovTPNJfzu5pyGOT5QwGIFsOauTASSy4UOb1JofCsw6V15ol1k+PJCmkCVfqAby6
NdZ834x9wwt08bbPVVa6j0m91HmPMSJ6YkypDuNFCpRwgcHzKQvGhakCalZBvY2cL2xxCHU0bnjh
M044AtDO1+++8ayL0AZzQMYoJmu7lxS2e+Rb2mVx/DHLFPWxArotKgTmK0w/YMhnK4J841R0eAYj
8siRST/5Lh+2q4vx86DkxhZZn/7yRv4kKjbH5tjfRi4J9kEyZoGN9aZDj+nemNP7cLwuxUfcnRab
/HeXM0XieJJm0vOKwBViPGiH9TupB/NuA0Wp50hsj0duJELMz5lV8eGcOvGAWXV2sy7abFOP5yDF
gVk7Wi4AR+8gCukR9/e2/7HJ68Rb0HT2tPY/Ql4HtxN2KCu4f6aIdXc8T9RYAaiMpA5V0rN6KSuo
FlsdPJ2phjv3DNA97PKiM1r9jc9Glsf0ETCHD2XcsrHdXhfV/4QPyP4BvdTIqcEc8NAeVgrLgxEg
ThFhZQFLvArpj2+C/bKrhsnDLDdgg36DzQHe2Zj1aQ4kcxZwBuf3QrbPVIhxx/7RL7L/0zfUoeXP
h0CMzIPQf5xk8e8mBfDCrURIwftyH5M0pjX9rpU5uJLHa3y5IHf8oEDRATtMiHpplUJSuKk4ALsH
zkx7VxAfuyNGZxp7D209lEGE4DM7tLt1HUp+gHA1Sz2AOsYuR32PC3Jak0SjedGllljFLppotmcb
odG5BYg5QlRb87X4MLVwMoZdh36TTUqUbzLhZCGGiEVtrbuMcZZkiuWiIYSX5IQVd8iDCXdf2KAP
RP2YBxK4X4/PSG4CJ8+WOwz9Bfnv9q7gLBU2VeOGf7XsO7C8X+BlLncXnu0s+LfSV771+ut7QEm/
qyFn1dsya7Za2v1k9bmvnltZqAuB9EIJ1+G8uyuly1DbyngOQ3BM35kP3eVV0IkozP05OahKmyF/
aE7r4M0T8fgcKtLtmVUvDKEy1aKGftF4nhF1THL56P1XMoa0gyzwNcLGCer21pCPjrzesxPk09ap
591ifIBLWmuNF5PRM0so/qzHBWQzeOAFW3ULYIxyCm84NoIr7Oufv6cQg5HRxIV1+6Inpg9ZYh3h
onjjbb5A+SNNf1dfUrfRqc3DCHm45Vojs9HYCcKjjmIntAfcY/4JE1nwaxflzC+48pVWed1AZY+N
ko/ry815jaPOuU8teF7cZaAUeuN+GFT/p0Ehs1kcVFSYyKTlAuRzFbA10tA00I6oxbhcFznHT3W6
tPJN3tjzy7/UhpmZSsk9NfVmgDnYQHNZ/yvTMQK69Du/eTUnox4bKngfOwD9BZliENtK5RoGXqzJ
E9rnA3Q71/GbzGNgyQfJS2xvgmLiox1qotH4Db/T+ox8/qvI91yOomGqNJMyVk766qD7hDoffDAh
aNpftn0zYPikv1mhqJ/YjkFsTR1N67AL9wCXOZIAkXIHLkJF7C3nLwVbfG7g28qlpSJIVK9DJEFd
oJIUfUjF2yXzNHn4D1K3cAaCIVTljWvBB2MpKTdt06QXDApEcMrhu7uos+Z8UQb0/IvKV8uI0ueg
14RWM0SQYlyl0l6Uzp5qGdJoXOCOI4OI9PglpyQSo5QN4Azq5Ad3vCUhFIpVxREpAcETGZ8+ij1z
HKhjKNDi8XHRAkFn0Xsd3Y5C0k2tJloy2bK+2kPgKdRkZ66bO7pXnkMmeSF3oyzTX37zDpAWgfb9
u9LMNSeL8fMz/PLqFmyy1eW0QU0PquYN6CCDMqebRTGqxPkVPcgdqgI6qI0f16sheSMlH2KIXZWp
W4goJEHpZrkchwPwwseKydQUnxxdeRwPV6Y6bSvcqzpahIy7WXUq8WO/LTvl5bmnHIWq99usO3CA
8l/jRcaYKrl6OJ3e87y7JG0qk2zTnY86Hb7FCHd3zdbBRCTld8avDHilKvDhNcJYeug3SCfBpwsh
uWogd1odd0iLh0O4I8HpdUXTYjpXorNG0I6UOsHakAeC0k8uH/xGa8FWWI1HGX8KJKHXgrnrXzlF
1So9vXier+0siYluywkybNnmMFZSwexiYDJRLAasCsa8q4E4LyVjRu6RBeqf+d5aqjUjty7u4eW1
SWWdwo8Gzs93TXrufDImT6wLJoL+tfC6Yb55rYlQ/8eqFjb0q9D1Iaj4lUzJxIPqU87V/Y2BS01Z
Xy8Dzay4KSYFoPt8gpINpKsjiZ74Hkqv//KPSKb5LOjiPFhdvkwWGbwl1I/u8tb75363sA0YPDka
/GfCsn4MQj9TrS3MIT6E49Ni9Nhzym1qfvsAQq7qXoZTpYwA8GeMpa1zB1dI9dL/OhZCBHAKziFM
+91hzKuV7DdY81syZ3HtUgJYNzoV4cr2ARE4KVLGM+FGynWBohXb4f+4r2rMOJO/pcEzT9MubE5t
NPvPywNgoINpGqCmcr3cObpKxU55ed2eaDX+wgfaQqn4L7mfLwInZswfUBJEnTclqaV+CwK2K6d5
EutaExTw3ZbLNdpbW4WLKoawBunuRALy1baDRn3lq9P1wawXPqpl+yjTPQBeBvUbOr43U0bFd+SZ
LwDhPRPgN2ZmqDoYUT2yHs9cR5B9HZqfwmqVqzORrRJYser3eit7CH9RZL4gYrLP1JsoxlsZmkmZ
Y7hDM3REDEmXPpJpH0Ykr5QWljiuwVmcaWwEsfQ8bXdyF5BCu8Zvpaak4MVD9PphmGA1nPN4XSFV
TqlY1zycbraiytUlVLfqxn+eoHxX0wFuRHjXB3llB+yjhmQA8UBpwZx8ZJUWr89hoaS7wo/m35S2
HXcMgEUXMRhVxMtCODvb2ZZ60KiwPx9RSoQPEwCYch11coxHpKJejjpAjbOAeLT7BEH8rkDZH2rb
LCN936W7Pyovmr9JcIiaFFx7wILvL2Sj+VhGBpueXidf8fNSRn3AHetQ7OKLGEbyV3iT7UrD3526
bIOLh+ZKJMHfJn/OvYH/CcrNWRVXh6HaGwtNSP/kW2zQj/xdzfrQRKjQdyT9BJgK6vu6mAfA4lHd
2uufp5PMfHxGZuMkOMLhDqroFsN5HVXU50EmBtcRVHAriGRe+97r1paRmnIE0O8FHhKzF7UiX5Tj
djiugQv1BKAjcmupq1xDeK3imMLPGH2b78TUb7tMzBF6lUklQqSXQved9h2kQirDUadfU3TWs8wD
Xp3KcjdIUpNA/CYqR2OoUcDj/uLbxD63h1/hICjfp0mJG3mrYrri46gQMnqb9Z9TO+pjXCXb+20k
VHk/BVnv8NV+OPe1kTx7IT4XeOwEZ7EYL41VVG0hAhUa8OgqfUVixifPt3xUd0SZe2TsdmotzhM8
uXDmrkBsEQwPc4ApxfehrugZ+63NwwDlKS+LariypfjWKSP4mUEwHITlqPs2hnRwM+jjHchQhj/c
AL1ifbm5q4PE+kY5lMRNiExqN2yogWgEce+GB5kZOTe9Bon+SeeLnxZp45DVq1eK60spmYPjhFSk
9t3N/R+haR6LSOqZaITC9wUUIt/CLCVvzeBLEnfxY2XBS8f9p03My5p/ELuNDLRN0ScKNiDD+JRO
p9ufWcuh6oSuDlnF2Bu8AFMLUOcWOkbEhO2cLltLf6hP3XotWc0fB5gL+oarU7NVaWHf6nkpVwfe
K16FKQigUd6CoyVjG/Ab+i0so32PATwLy0njeenC0FHZVCQu96GbyYSbZhSOecUjNHj2csUkxkXA
2qfd8vyhz3B4i96fJ3ckcvURQvHxQ39XvFxNqWEwfCxdRLlJGDi2Kfcek3JEah+3uUUmY3p4jXSR
6MwfNQgpJXn4Jxi446XMI9oPTjNmmG5dBMUjJT488Zm0qD3Rhk7xLoIvBJnnOLFU5P9yLHRjeJ4a
KnB3aWEfzeIoltqKnYqrRbGwLGwGJ5QFqMF4wByWRwxlUsXN83ckHIaLW8K1F53Zd+SGGjmHcvFH
2zRSK0YsUY8bJCx6+SCeB8qohwNsuBGpPAHRcRDUbxptKXhGzHFIG/o78StfJg9JYME810QXk2Dt
EoQqljaKlewWHBJpdoJEsJJa4YaUSCuH7cKwF9hTCCDtsU0VOOupvNJFcd7+why+PW15Mgr1E+lW
OZX2a1IBbElRXY5B7hEWdtzg6/dmTqNgDoH+bEIbGFXHxRlbq7PD9u8fA8/PNFE+3sDPjLZasCJ7
TVaW90IPPTvZR57s8hHRoTLj88bR7xXxRNL2IAAQ4W3xFPLY7nsCfYM/OX1k31eUlugBvW643Tw9
YIWLacnmFxLJcg9mCLWuGO9HUkJIpOJpTFhSyaqjssiA4Hkrz8gneFrhD4HEZEDv08q6BrZyG0OR
W4tKGnRtLJf7zZssRCEjdhw1jBjWTYSAosPudLxTsh9gFWrvo4uuSxlng6aFYSE6THBhQ3ZIzwrv
VWZKbHeb3ElYizbIkaWm4UbIXtkoCaEmKJWkNlzDcOF+lHzZUeFMjKMKI02a7IyiiU3VuW2sfmEe
SzQSpvKcAGZcHTOsu1f9XChDpG08VdYLe2ODaGyMH9Qa/ePVXnT9Tk+RV/vG48YFJBhORqduOH8Y
tsZ9Sub56TQ5sIxPNvjeNfUVBT7874wy/ghdYr1p+wqIiZ21fGCutSGjbaDHjecLNhW3nqltj5R+
p4ACbT5puLZS9jqkVRzylukGSxQcu7M1tOneOBd/45TMarEjt5kG6pD/1en8K+S5NYnVAr0FtX+U
gTfTUu4mTUBtC+MrsWOG6MpC6RFzvL6LNhiIrAejC04CXJXALWjrbBXdctG2VCW0yiOW67bJmWTq
gtTKi23P1VEXloSpmgZzFv6s+K/ElNcvwxt/dKjotzAftH4bfjeuB9USk8SaTK72/fQZOO13Iaay
fwTZRjqZ1+zHOAYN1dUvV6dEuM6fnPWN79o8nb5iqLBu6k4ZJ4sjlaKzJ0gBaX4mG7PQ6lqKC+tI
/Xl60v5EtLhP4dCYhUyCewalE9ARTPuiYNzsfPSUZrm1RK658JzI+TPjVC65qiqO/bmmcQ8QCIT/
cql12z5gq9VqCRl6A8GpNpzTIKPdv6bbJBEyo4jpL5OCS0HZhsDdk0lfgHn05UkcY5SRhERKm90I
Y4UNAzZSqUMjkWQ3XoFuqkDWjPhWPeL5YCYGJGKFRCOK+Zjx6Vhtmt+MpqJI7kw9/FYmB3+n6i2Z
lfUAe4U3Rfstnw9tKq4kT5cfuO3CZ9qbUYMAAf9AvmuLSKNOYK99dQ52/C5SZj7N/+lRU91UVp5E
NajmyOWPRdFPVxbzXJDhmu2xYkYMir8PD/SuLVaNtQ2YbK847IsI5iDaMiMhJnKCwBP6/KDAjYWE
kAVXex1jGybWzYXEu35fOQA3UauZ4iOq62fYfzB2Cepvzlz+FDHhADF6l9fK8fD+cmkuhsLJLoPy
y3J86G/n/sIbU1SC3M8cwloviFN2ZEfxCMALbB4wowHu1XeWgndQhI96KIDTaLrAP+dbJ0CFBpSS
O1aFCAhJ9x0HFDVfjPM/2UUaDSkE5xPmPp3JbbrSCT3vmKUubNbjFFH2ZbAf7V9jeOhNZPSKG52B
4r1Nyi7z16YGTDGuEM/51a9Orfz+sVbs58bpADoMXyG0extMgzCdRQYhUpETpQJCp/stCwYx/2Q3
CLfCrSk+TP+Mcbc2oySv+F0cl6kcA2+tw86ADTg6jNI6JbmQplHbH07dhpN2ePIWISlSNTFq6Rs9
setjUQ/7kNky9dXr8iKYKzZizRzgRir0ciRX+nX7+QdHukYuLsw+Etsljn70CkLMrLOskfJGaAnN
J6fTOYnK/M+kqRE8sKmmoL2vE7NMNW4OFJ/d2tOGm+Y4UtFBk3MW06kJO0WGokC3COwRxU0nH290
jRgC3ow26xV2Kyh4SBJqtDs4tRxp3FM1Er1xjbvJ1dMIfbpgTTWLpyqF5knjeCm03K2N/NXIN7LK
YvS6zcsaHK4ZPaMGzKIUs7THcziZkMza+TRtgrxQlDFqowV8uEqEpJD9XHOOBNklkCQuafuZVVah
H3ZyucQcW6IpCMEQibQBKpkF1n9h9/nxdmsL4vdagEk678gLYC5DyxwW5CflOvwoSZsLsyCKvIiO
stIxMwqL5tNKLoJvA9PeiBCapR/JLeyDgIo3f9kJj6zNS2kBX4P2q0BWsQDSK8c1n23zobkIZM8T
QFufy92b3hp3e5HjOIWEOhBB2iC0zfq/ZUHR729RK71uHMhL08nRpBGM4xT03eoOTFvPgP3cdq/H
G6ym4TFKLdkfcPIKq0ONuOV0947/YOIzBz+Orvd/uoabu6WPJ33g3JKwnfAQuoHwVWnAKh6aA5jr
oXlqfKumw050xUkXVf7ZGPloNJpd79uI+IKH0KZ7yZHwD3vZMAL/7rvZUH1+cO8Yl4QE22SDUtsN
MAak8lysH2BwEMOKDT+ytLOfEGnzehEQN8tVT2hU/xSMxZZ8vwLKR4MJEVlSmNzPThFn4vMr8FE6
SZjBX2cFBPVQl1KUrPE4pH6NeL3jr4TiQYOvK4bTF7+dxlTBKCsZ2KDOHhxgRVFVp9gtkVfD4+nw
Dt98HCekE552VoIYmx9TZpi+l3KfQWGXN7eI+JHsswCrbLxsMAlKBab+za58GK0T9gd9L274l2GC
RDwvefNtteyt+ksUnA6DDQOT2bs0/3N3eZLSKqEN+l40+VuoJP0XUwCdmsXVZnUJwz+/rJe3APxU
jbRVRc/Wh3VnwZCF4EjsXsBjqFu4bFplgxFtreAkTCtX/C/KS/N5k4Sf/uc39zeDnDz5m//IPO+q
Rn+wD+IOHe7s3ITC0Y0obKNjkFP0IkA3dyCAU3GqGxTEEsHgpjsmsfcD+N9xcMbfRPfeadtpVBS3
Xx1aXWbhX8AkOcjUz+EH5yjP2t0LZH9/lN2UJTnp5D+IyPMDCinxju0G+r7wfMBhUD8Bx4xafMf/
O7R30iXm8WVpCQmC9Dtpl5OpGhnB2S2Wnbp7VmzqA4ED+JXLG3YsM1RS5OSa7c5ACUxuA9DLUe30
BYsYsTIMU/Z8q236R47cHGTkwfUPugglu8FAelVhm6NKp0KuIxFixrJuj0X0KuI4PpmbVz59kfsL
NquiVQFkgUum/07UC+89wzhaDKxWiBmDWkiKR1fTM2+A5y3cQv840+juKGvE6iRacz2cZUg4CA6g
flKVTR7almmGtJMP5pJIxmBPlt/jIv3Oz04gD7KK6bYIB4VhGECrwjVvEcVUENmuFhFOCn2J+Qao
YGFOgPojSvfWzgXUIXiIjGOGFdRcpbpWlJm5q5n4OnAcAKnwhN+n64gZwReQZEtDVQx7HIHe0hWN
R7vwNQh558xDVibozKJskm9cUBmFTvu4XyyvJGkIq1FiP3ZjtGbYoMtatSP+VAXg7DMTHR6mz0+6
m44Tmc3Co4KrkJgNiDg+HbhqJYQhrn7jilxflu8BhqKVgAR4sWygEKqF5HO44pg9LPlxxrGAFkge
h/ddPSS1euU9q5t2VHqfzfE+jfWvxWP0T1zdXmyOiIL9BNp2/DfuIDwxIodnmO4HIDX06nF3AL9r
oWa6JL97ZzxISghMhfUPoVOA19T44dbffLkTo/uBiKVuaLfOS8pMIpVJFeBz0FupZZKQgb2OZa3L
gdAOkZemPqNRBLV6AK16cKpUnWMwt8QMaimJS48IaZsYwxTVRKr3W9683/+3Ki0PRme1cMVZ/Ilb
ci6NkEBSbut1o4VKSfKWhkRvplr8Fayzkl/XKGiwxxHGqrGMFVuYhlLrW7H9nbuaW9ceQqE46FU+
WOKuqjUczjZF85qeuCE4cuNwifCkal/eGo/CUlI8/Dt1dSH5OQRZR1LGUX3yB2KP6uvUx3Q6hUaw
V0t41D9c4C9BW7HIKRuiibg/+eoQha3ip81JQA8yg4S/h5xGDzt3qQPV+/U9lDdclurvGP3EmEPO
XboM5nWEMzrpwHa3X5AdAiRKNt/wiirh2Uu4WxXDPwmdjRr8BW39hOzWsgRRFcXzoFv9hSbyVIzv
DI9UPZBb5wlRqHWVKTwuAUFNsut37598/oRubmWn02cM/GmAvnw7A48YZT4pCyONVmz7K6xB8kE8
hfbXphNXp8q2laK+gT706eD2Kmmnp70idpbp8qfl/vtEjUzk34oMFECyY2NCjaT+KwqgOiQKUNyp
CK/yL3qoNw20R/193GRDCztq6BB4IyG67Lmjbx3yp4QjG3cP2JZ0+RKY7z/HwXHiVdwe/Zdf8n4y
hmIw9Vh9ZD0J6vZzbTptRVpD2d5NpE1N0t657t3sYI2dqnSpDAswPgcyOwQmQAapYcQ/dxpKZMu/
gp2gu1mS4OGnFisyWclCgWOXlXxQiJP4MA8TN7XviztS3Vb2a7prsMeOVo/AzderorZ/y5Oz0RMR
mddzyH28jCQe44nKdE2j0k/01RpKF35de9vuYPz2uZqS73gaiS/L9zwT2ZgXf6Q4PTZfSPQEqbFj
EaYlGVPs9mMWNMikuHxAP8qccL5YSznsfSOu713l988llib8ORxAkH2rNrpvUBh44MeITqobcgfX
AoBn/bTn2EBVlxBNu4D1IWdhpyRfwtDz1pP8NpfcxaAzYvvFuD3c+ot0x7WTmd/5m7mmHx1hbh+I
wkefBfZCH2YLPJd2qCtmzrp9qOCIFwViqAYEScNhgbbBpgH83utziY/P+WkkJr8iQEjfYu1ebBwI
/htsX7np1WNfkuTTv4YZYd2ZXiyFwq6gCBLapacjPtj3s9tCDJhHVcvyGtJv9Daet7OYCE0R9/GS
+A3VPXP7580j+bYf5xlLdnwvam5BBhe5GbeIyLjH1Ck62wFrysDigsH1GW5/k8QpUXkH+1SM2iTx
F8rospXsSiWETqvJxTYDS9K6uEK3tnAxJ4upTZ0UVCr/Ml5yAIjjm6CMHd3TLpU/9CFp7jv2MLiO
NBrOI93mUmo5bm8NGfSj6n/sDGpARBrB728Fv871RkLp94ASLSSV0PnI1dfnpFJQqlwMuxXLq9w7
GKt/OB7uSFBB4i6GWhUN32bK4/toPRSFw7R8+SaCqjlyRL0X06pJbfI6p23Q3IkhVfDYAF8h4abI
wkolLRRWYb+Dvk9Oo4N+vwPwpuBX3hG5VPr2sG05XDvFyLg48vXdM932k0iSeUGBtm6R3xwOgD4Z
mJadcT/atTrFbdBQl8tDXUPzZ1bjnyAPMHwHT0iC7Iv/YXLv+9uofV/bKzTlRDOxDrHPGiD91F28
+a6bPrFjFfLb1KHlEVcXr0ypKC1wvBuYA8lcxYT8uqb8U4MpfTfyZyDZ5xb9aPneewk9398ZWD72
bF7AixPUM4s0/MUhl/ZJ3ZVAGJlW/Zve+sHAJ+2j6mAc9cHp9itq2YqNxEoLlQUZi20td/CAEjL6
74ryoNsQxC8tPlE/xa4UNoi2DAeofE9n63E5GHb1KYAqRaNfPGXqGyx3veyBG00LoPHRayQ9wDLB
TawHrpaFL5n9I5wsP5bUWMOHVvIhbw4eS2mygPEADQcaoh58oQz5sk6b5e/lRHu9Yh3HbiX6aSfR
DAyjvZmRbilvrEVRXMGd8GqZJfdS8EX76NxrI+FqMBHfj5QCZ83EuWuMbWcqoT8z0Lz3dZFfvet8
OyibVHnoQlvEbaT5ZA2uIrYBb24NZ0VQ2iimFHI9eyoso+DCPXvceidQOfTJwoZKrKbV+2N/3HRN
Y3wws7sK+FlluUL0OkJ83CXqBG8aEUY24DEWzwQOrrj+IJs7AhKLLwfobThsQQF7walH73QzA92s
mseE57fqrnFw5KjqJq6zZxaqOwfxB+CY08TAY3+rmaBpZtEX8s/S9eHie7xqqZDMgESHNqcIY7tP
KdFbF2vy3QrLg0EUk1K+Evn/Fw5pEDIYWDfXdITmu8PrTqqOBjw0hhzU1TC3qqhRV2eq7WygVVpF
aQiC3/RVLZrvmRqU1qov+1dAGksj8M/0xsJqEOXHahuXXWuGoYhi9hZ5bxGNNrh6R1vgTweKNIGc
ymaKsvLZffhrfXyxu1NRBtXpjNLujqJVxTuxJqdAjMNSSrcDpRLe/fZEB4p/loFtOURTrg8xd4Jp
kdMpSveMFWYWDdhkwOw8fl/Yz/kTbptQLWDLc3dmJfZMf+eCJn5JmxYX4ZYUKVMXxFDT4/gQ1xJs
m5SwbNAjFeWF3qiVtmE0VpYOY/ttGN2KhCPix4i9t+EXB9YLLxhv/7cy3KAPPW12qU64llDafOzf
uWYg83FLH77KB6OHgiAm/ZUDbNX1vKxUOpuGRRYcp5IUQGnkLyriKSqfO+8fJ9NFLlhGuAUIhs/N
KxFLoTRgvNmNnUzeCrDewgqVEc5JzvTCuiP/7MffedRT649m2r44vvOnkM5bO5wWTTPMDElxn54F
R+y4kK64L/dqPqQD3KcWx8mv8iuxMgxwqNhLnYmBTiIhThFXnvmvb1HutgmpoRttlMHxUa/KplYu
IuSCrOFHi2nN1Fav1GkD4MWAWBMufXt1NxBD0gRktEYYQ+FTjmlYcqNXlLCE+OuauHzuUxlJnIq2
4TBdWTdU26zABw9THH/9LlCmjTUb3go4JwiDliOdfd+AEs4BgZ3Epq0IaJEDXXV6QPM0XOhfMrEa
CR3MCCrb1nW+l1cKg9UMZyxOnN921CiDY//qjf6nv6WkO5QAxd9b2/MtNNkWAw7PCta0IThhbycY
sLSK1G98KmxOI/mGgqFVIbh93+0zxMfjc4OXLjzA1Q/1QC8Ci3dwEOEWOqyO2e76Po+r7S2p+KvJ
c0nqkXUr7AuR3/MA95SjdlobyTdYpBrabJD9yn1CDXdhPszyBoruNlhHTd7WcnFphxdfBOh2dzjs
0tPrc5sx8+sJbFmdVl01aqS2RTA98Kz+oHRzc+pF8u9Y1oavS0Hn/rgpM/Ma9tjIFl107gKRhNHy
5nnLZLKIftTz5b/IeKS57081PnTkjtmfbJfsspQawYCsnXc6h5qhp8vH/jrWB6gIkxfAQZRNmolf
nAhgNfyXBH96pzTmFdGG/WO06Qti6VMTTTUu6qdjALTZGw9l7tSee9o4Mg0uBlq10pRXmEEycDVF
u1vLU2uu7s+9LsDwFpZain34sXOFgmveQQJGkcw0B4SZqimplWfPlvwlMHBSbeU4SKz5miPZAgLg
bLKKVssgzns49s23YpYY4w0ve8071G6BGP50XIr/bH/ZPRFVx3lpSTODCjEp2fmMiCRN6TQ5+gIX
Q+5YrVxmXbaLzaCWeeW4yBtUX9Rv75CnzMGfqky1D5f6QvM7d1dHpsRR1jC8GsN7zP027aPG3s0O
HbdeFcV3OZreXhO6a5TfZxuEuVgE3JZhi49wew/A+09LcVGJXpSSXCPtZNPgKcGxnEDWcP6zIf7u
gk0HSrNBtgdP20fLXMHRE+zItEc5o/gMwMUIHaMBgAx2SPvYN2Teeyb9dT7FUXhuoB0vajBoSnGJ
cCXyMIga813v+5cCppDqBLn94XS8CuiufOC+MNZUD19j04gAlO8jjBndMZ2UBKHTsaAAhuiCATdO
80TOLBZYgWPGjBcoJL5Wnsku1TsLmPHVNIbh63f4mFHmwRSBs0rmzx6tGx877cy2FXfVJr1kmT6j
BOOoLv8pb0OANc0s94jh1pJghZWmHhponHDyZud8Lslhq15xtsdPMii9kTKhwcYml0DXUcKgXOOY
M8Zq1WGhS3NzK4T5Ekh382S25GK60fRD+xDKyssN/JTwrw9oEwkJ0PhCq7I1HyZ6EGwgn8MDQTe1
+LZPGn8plUbmfNzF2dhMMMk+2F9C+Ul+O07WsaITSFXIeig6S7RCtn3yZdg6eRJQmLx6AIBpXnDT
SwOnC/7CC1Arf5Xri8QxacoRxtJ2qitm3VEMLGSy7yqu+GlzYfKdnbigJ1wyX93skNWtouUwz02Q
gzRfldujVfHBdVofve2rOu4R0fUXgocK7kPAcXOb4iiOx4WPJH7fgbSeWOFSwWzDp8hSTkBOhG6b
c0OX7yzhhfOZ0BkyjrGclALYKnGbmcwyNycAQ9gGmnopvma1wmGzSgsdz6wCr5X60oNacTsTHdj3
27ak8l3loF+Yl/Ava3nrNkXwS1Ux91qpBw698bmvtimVpm+csreR7XVRNZ74b44W5ohVoRkbUAO0
ByG008NFsqoWdQ7gRGIFMDo7hw50vtzS/S5y5g6SeGw2vXUdIC9eEN7/Z5ieCgBj0OMXsORIuvq4
CqMGR7CKCZY/kHNOAolo3mTi7deDSUyn8rBrdIeFFOLfETeeMiYpKsQNgOS/99cmQeEFAD0M88Fp
/5fnm7FWEhAGC9NrAYKJDPWarGNqG+j/1+6NZAreUJWpUZM4eEOSZDjpZlJkhV3B/THm4qfFl/ij
4dQkYJ5vZtvKTYSBqD1yoOl1GiCv5LiJvze86OaMApGsLqnVIcL9/q5l+z/8N0QTwwOphfp8wup4
6U4clSRVWYwP2qxJrk7k/vNDAA6f4cHD4zmQddUYiih7m7jON9MsS0KjHI1RkCK6Sfe7u2lrdhkg
MHEoPnXkao6KrOBmde+ogxhFQnfjI9s4i3sGs48CgoCrSL2oq24B3Xl8JFbQ0t8ozbORhUGFl0HX
1EQfPU8KCgpFRYlOibVhtP+LFVzsF1+PgSVFWpr+W13AsQSn8TYp97J4wX3yHgQo7koGJEupBrh3
fMuzqrK6UmNSKK8Ctb668N/Rtjr3sWIiAc3GvsDnKERxlt/ICNzEUGdfIm982YGnxolCdYJhhxPR
tHMrPtftEsoAo3SlaEZ2mW9wsK5gNpDiSJoozhD0jLN92lRqf9l/nQRcV8fRZm1JxISaFmVgk8P+
FYPRB4sbYElQVrSVWQilg92uRm7+Dzlrft1amiOJvGUgYOivvs7eCZQ9Ff9rQZzQ+sHHi5DCaEsK
vaybSStowJzQvhX4IJl7EZfxtnoRcOoZVXmGbfgq3IbK1vMnNvq77WdmaW5gvGwL+LQC/8c+MBCy
NAbfNF1Qy5Njgw82WRQvmfbyG+NnbASx0QEL37o5W+M1mXeOOlHVWGPqH8lv0Ex7OSDB4VGBEOcu
eEYVYEJGCUvYxe441e7+kwxbVBSbHHXXz9kbQvcplS83d/qEhCC4feE4FHZTIt74iE6/TCAX8RSc
EaCxz/VFom+s0VpNoSdwvvqglmW3q19UJRS42+G8a6zRE6tDF5e97CEmE+1XmZuil5syS7QG/zpU
unL9+z9eg8vc7FhRZQMxw2KQx0ealgOg2E68s3sPv7DKp1r5SvxXCHy6TsII+PGvy8YSzwf+vxDS
/dNy1MtI+vMFnsKiPokCyAckqL/pINwHT3xXWfuFSJawX2m83vd3ifyZQ7yt9Gx6GV80MysaU1ot
44alFPRNoKUVceNTT3BOhoATCqQ/wVE15Fe7uawd7t6G2KxkfvUwGq5nRlgr+as/fTupOe4dE13R
qJs+XEE5UDvchgICpoaimm/cMS44puPhndGomGDT6O8EwIRqLpzhqaqerj6g+Ea+gvEMyVBnxieB
xhvAQxZrGPYe3bPlBxqYD/NwenlBTxPikllTG49v+SRZ6Z3mAtqiXEUPL/IIqloGY78FdMUi+t+S
j0f3gY0z+dl9OJLWrh5EaabrmzgFt8XUS1hsisdw4Or8zaVm0mboHE4mPgMilqwKo7Yz+axIPu1d
ObJQbCgySwKknnrwMiCSFPi8DNloR9+nycLpCTU76FLwhmOLysrFnF0dKlzEuHvylCR5Y6ljpO9+
GrW+MyrBfh4Gd4adK5Li+4uV9XS4up7+UNCHCDlpEC6op2o0SqfS+Qacbp6T1Z4+eoAebQQ4IjUj
vOXZ5L/xChTRkLBfKOHQR81pB1eBFiNZNli6mEMcyFLHjpSQF4LVMM6Qk5gKctHfPnqZvU/KGOSP
PGf33cN5lYsL/VN4frihJJnFxk+Mv7RX55Z6E/UuVIGobaaI5BTM9qUqmgdzRxI0bdbyIq67JYq+
WS3qrNOeLncJtx3S71utPR7jLIclYbIRu74sKrnQrhNZehh/4k/jr+UgrH+JHxJcFFCg7glkJzGS
khBZbGL4M4X/d0fvvoW2VB6v4aRQwrE+PGtDCUVoV6uO8vzDRx0MACEuKJ1O4h+kXX6ryOQf+Pim
MB0xvaHVaIoIXi17k0bay0BYakHn9o/2eUcItSUZHD+Apd0o5w8zLRKd9VmB8iUizsFxq4Sa+0+2
ilTTApFi2f+z/AtGQtfRJkY+HlHjyI/48+a/vTCmb+6nxbPjdcZBTBX5DtBhh4QejvbADDcEfT1X
n1mDipqGsZbPw15JNEwn34H68q1rxrdpbfKe4MRqIE7GMzbQaXY9su0IvijI9B67MV5ijX/fcCI0
kRU0L3PlM/qB15FCHj3mI8/Oji0CrMm/O0DmjWZNKa56rOd4ej/3/7Y4IDuCEOvzjzeEG06MB5Qv
RQ0nLyldoxgPscfvLyoQumNiYUob9BM5c76v9r3pOTRfM+UfTvJ+K5ja/UHfWU0Brgo3/5vQK3/h
UJ4IvtrrgJU2Aol5PuCi+2+huXswZ7byfXwZ/4tuRRKx/k/sBnMM1rCleWsa9c5cAuRYLwZskDDj
6ei+fa7Qz2X/NRJ1TJM25bTfxRTke5i56XCcbpKAWDIe6I35nABCWFL+UWi8eR+GxasqWJU4JgIo
5tkMmT5hDcBMWF8LXuNctYGhufzb4W6+y7TYL5PYfOlLSpDj2HY9X55K7VB75EkKT/WjJlMQuECr
FhEFuazxrUwzDkRgB9FNtF8gQqXd1PcNSjTIa3TIvc4aj3pLCNw5c/JLmc3RVdlejeWH/fgLk94a
utEUVze8zTW3mcVjEJq0c0eAPADKnUH0ZDNgtR14HjN8ql7Gd/gEeKXn4VSUk35EMPK6Ett7s065
sCp9V9zsPqoBygew31160rW2LOBIkKZCwVkpFXtpCNX8VJx2iOlWJPORnK+K7vyMgtssI5t1DCUK
t91TRv7K7GBCkTNh21KB2m2L93+jFeck9J1A5ouu/tGjPXlGAh4SoMFRMRsKFqx4FS7zhBgrnHS7
cGM0m0imMHfgaPpqd2VTg4cGhn3PWuDTQMPiH0NRRz+mNfU39Q5ITYRILUQexW6u3JAQIPdyzrJA
+QM+nLE2qq5NP4hS+yOTwodrGOEhOh0KZEDmPw/fPrcOUaTqOZNEexNhOoil1siQuoOh92K9c3d/
6lO6vxUSfuOsLzNYiMZB4TfGGXVoK2R7oe7PHCrS0ucmVGKal1yG86S1TL5PqY8zV4UeixO8NyH8
ijhvq1frDsH4heDoyYEKE43IOLvEtIQ88nQXD6Yu2QEfddYuaWRViTzOK8JDmA43aZP0dIRgKTsz
sPe1TP1NnfWQZaRs07Z4ZSQv2hbfw6qhh1uxosf2Zd7ll6ByKg+D0vW3dtiaLjIbTNZwsBM2T+Qj
TEgYieDBMYXBelODw6HHjjL8algPOoy83ZIHQ1yzGuCCiLSB5Ik4KSQq6VDAwWmVxLWEgEuV8Qnx
ykgzy8+NPLVNLdjBoGVpjn9Hd6QdWn7Cez1W4w2tVo10qWBj6QUnazd7VbYPWsSfA/hAgR09Uy5Q
pBboxWmHyb2QOFudgW0r9pL2HXdhJDkgxHxBj5nkVL8bIq4QZnZIzix5afJh1Y6hscvBYlPhFEFV
oIoNKFTupPKtXa1Xqd9Hz9K8+ZCrpDX1leHkfKndOdCEKKUzYZsZXKx/hk4Cm83A7aKx7UbIUK/t
BoWMFcyZ759QP4ro8r4AZv6gAj6AbZfd+D21KrGI61kQL3uTy0SBrbfrDRbMBUDWdTl3w3JGuUMU
pDePsRQlvPK580w9xR82wNTqNxnDUwCINHTksCM53UBzKkWjYxUkY30Ou6vH0BkC4x8/E8vWlfbb
/vK9CRf/lm4zYspL6L3olaP6J8FZlpp8nIx7Nw9vhDlUAtZ7hxrfjVj5Pnh9zWZdIsg9Od3S7fLT
ZLH5eliyN5dQpAk41JAyvKLD+4gOOR9m7nnkdfQXKEEp9/DD+HmUEjkYBKH7EgaSCVkMmNZmh7m4
c9zvhft0+K0K3HSg0Vyq+F5riDVQttVXMkk22STknC2RKMBIA5OSA3ydRZkfwlQ0tdYQoBZQstt5
9mqGRBnSU6L+ed6iL6qAFK8vDa3rADajvZutTH2ggQwT907RxPbcBqPdg5/yvmHs32fLPTU/DpGS
NWH7RuuPZ3zf/mwBXV9u/lzu366ipC7l4/rPE3wvjWUw51UuNjMt7Nd/9t39DNChLzscVhPr2NOH
ZHjvsYDZzi3fxfkhbzPaWeQWHUhhTOdaNZi8SI7x0dFleXwiankINo2sEO/53zHF90e+Dtc5Uil3
A5wf9iXblBb9MvmEmQhz1GohioMNHF3Q7D5Lqv7dfxP/qApZAagbHjzR1zaceD7UmMwnzXC0rKlC
IBZAaXH07y6oZr5N1nYjgxNhQrCy5BjnZIHcqX8nqCpjuZ1PadEagAUqrJQAqRTlruuQ0r0lAUCD
uLpW+ARzP1XGCVfFpgufQIcz4jLAsMfmBWv/3Rgt3vf2f4DNZJOqStKIRcULaxfFPfHgBScOqsU8
KKgmd31xtHlq+h7avBegZuSO405OxekjhWd2lBydIsoMSP/N3Wb6F1mMerI3wyI6Vcoq966YiXHZ
ad6pwceUD2k9rlNc8No6+RGfUKp4QgTmvyYIC3qhMQwIKYq+TC0zeqMxzqXPkJaKPwE0VWRK+fN9
3rphv2llTzOIUfxoP2RS5knWaK4DI5fShP2d2jfX1b78h7zrQV2NtGRL+4PRtr/UM2jGy5O+bTkB
L9SGLkN0LmtQddlt1UNsM0FoaO51B+fO56o0t6Hk4mPdEgFDnTiS6UIB4UXAem5ULkaK+Sz8B/ov
dcrVndAj8Y9sOcwzaviTfnmTCKbEtTUPwwkysg9NxYfJSAlvOijjYQtqVKUVrNTIU3md00ACxKWc
HRuRiUGVBSo1hC+O5UOZR1u4fwrzRXprXZWl72NpY6bZ8bKVBRilC6QhN5mIUhsgwrj9sQ2DYgMF
6ySDS/pamyIY9PYO9DFWxOHf0Y/eEtQsTl95nxdK88lAXO6hgM/HiN9rDhgi9fUE7icDY0JJplmW
wTJ2OFk12jC47TXiwdsL9eW1hxea4hsOAcwwaxINwje0TPB+HAGr/nu8jvxs0RIH9vNux3zbnSv1
Zw9OYSpZy74MMN54+77TxEX24fCGVAFbItkSz8gBkERfmx6pwJZ6twzy3O8HaYq1ZhJ8GP0xP0B4
2KatKaBdGqwQraeT0m85n6ARdftadQP0xxeGeSDPCuaHKYeRuMBP15u+JRh4z+abptjRso1QEnwZ
FXJdJNMwLKCtD0FmMXLwZxd51YquMvD5xmCPceFFQc4NIUt2t+O/8DkXrywyu7EqvH9f4pdSQ3o4
/gPsaFErziAkXXfwT8Kje9tVAlA4NhkWi0wYMEwae6j6lXKSLDBCfM1syFE8FBtVgKxz94JsVkU/
yjN0CXC6atSRsEOgrnvHx8AiX6zKNmpmdo1/XDYDVW2vPv/bAdzEoBwabXHlTiv35THwm+/3ZTtz
y72UBEqxgWbXLhWYW4oeeqhlxaBOfI/nzu18WuX5gTVjF4gJluUfu4t4idF/f25voH9h/y5lH70f
OTqUPZvqgJKgb9GpuRcN16pM1jUrzALph/oWCTXCGb3DMAKdrkp9Hi47fSUd5GyIVmk9HcRHeVQm
k5QEkY2vI9OZxNh441iCSaaJmMJnNntd3ETdHtQdt/+cENxMUsEOvvezD4UsrHtmh7I4b0hydEuW
ZqI0wWG7zHPxIHUiQ+m5hXCBLAa3/27hVApcZUZKDbGDRoLte+Vzr00C5rHLlbW7vypUO7a3eHWi
ck2kxN+HM66gBn96HvP2NUl20bc+PEGr295mvfOqFxkfmBY8nxmbD0YHzEPbeRBVSf24fb1Es4ye
D1VH4h2ckS/bDB1BPbo/djErE7yKbF/LQ6MM+O5F780E5Aw5FSQXEGu2+ClA0Pj55Cumssb8R4Ib
FTUN/j3PrBy58Ekrw/ySNr9Wg0D0N1srkrvjku8yNPHBpsM5jEMEmHYSxlasbXS/2rSWskE1pD8+
NHe/tzalhD8oQM6c20wbBCrWo4MVmM/j/2c99WIR12vUGf3aiAzF/UsGJglMhtMMKRsPlyNE7rF3
po/uppDV5aWzjUfrHmGZmrHXW/jnTVaQFdJcnD9Dez4teKmqGGrfHcmR61ewqB2aAWTz9sDC1C/g
aH5BT33q92W8YQ4RGs+HvGa9MjyVgDBsXnTxDen1TV2PKYfLlHvzbxANU23ZzhSPyQVhuLgh+nKT
iyM2yTY6Dm/3R+1y9+IDahR1bAc10NdgskXyaMbObf3tHIxZQFHbXimFYklk6EzB5+M9bD7R7fcs
nwLYwmSPp3KbYWPCCoyv2JKaAD5KfIqooLYny6GSAM6txEo7UQ3cmRNkuwdE2hlKUK7K4RCWAsP6
tMQXce7PS5wvCIxX/MNrk4UosKrIXoo3cJFzozu3B2NAcJz3CiP6GhHPoazHcRUKDSaKa/bxMJfz
hJZ9x3C03CDR14ktBxZsqv+HVArVaRH9gUF9HliBJPLSIgah7tHbS6JBXIeTpaEua07+zXRDNay9
4p8M6bpBST1dpBJgSnJmmBOwXEXj59zTi4zmXkq5p61PWNrxSnFckhuwsAnSHYxxIPMu8B2Ijrh7
99yAzCgdIx0aBuX5+VWYss190OmekKwgQp2BIE8tGlcy+RSAkEW2Q1YPR3MkUgsM8pnkVVD1nYWb
lB0kzXdPQPIoVIxW4Q2wDCin0a6hS0MtYqV3Md+Tn3AR4+/TU8dYBf0Yv6QpV6tBeC9snT0/d1IO
GAV1duVEo5Q83m13DEm4JyH2abDTHgKzG0NUfLoNnpZfkk9kfvANQWIZDSsuOIF9HuIzYN4vSiWY
j7h7Jtkz/ig25dBUikkWb6zlcy/pz+/8lu1+Mte7g/+DV+PEL692HoQMu2FylbDF6k5/zTrjbfW7
p/CZ/TecNoz2pJfK49m2YhHWeYriQVb3KhNd7lC8/R87fuXB7Wn86B3v4x+ug95Vc3doubNqMB5b
Nt99mdw9kDe/uanY1mlFjVjC9B9HhqX/KK7712SgNUmWrvqKsWBhOV6YcmnNQGciEKA/ItCFB6vv
VYHciiqqPmRsgvYUw/SrGI+lQ9vkq0Q0MdC1CxiIcj55RnMS/tDiTWWJDWcYY+3ODlfW7iIKQdnP
tSzR8VxlFE8am+Ys17lwsfrqmUpx/1JDDDt75M1zNnUkuuQf5jorL6hgCFAZyVyhw+vRsfxhaawJ
8x9vhMlSNr64U5aXr2vVQ9I8D/ZxROg2tfz9WATR0tsLFI46Quo1KJOjfG91fmrWwN+K5xoODbi/
DotbV6xeB3tue+9hnjekcgmZ6n2wL/QHClH4L4F7ylBLOC03nseOw1/54iFtFM6XMQF+ldIgrHv0
WoUi63R/mj96VTUxtsCuBA8LaHFbHUqBbERrloK4IhcvOplrAxDBH9Vq/udTRrB4IKcTzRrYpPk0
lkXYLd1YTq+mAWF6VKSHVFJIIAOynmFAWGt+BuA58qIZ1TI+0M/X8kpCsu2spmKwHslmCyYbgSn+
Nd4C+t0kzZqSciWoJv8eeRt8GM366tmsVhxNgXWqRwqoFpxewKhgl61iqMIEtuAgyymdL2UAUfux
badKbqlnPT4jB3lZu35HZvMYVLmiaVd59kyMkvUIbLykyC1OdIGjknRkxrv6Dl009S8uLCH8jSne
pKk7El+mr+/fYZHEQPzvfahgpe3PaC7JByizJJnx7ac7YK/B+qyf12ywMKjImH9LO5T8Lt3tAakv
WyQrSgj1L1Rv1jBY5t9ya4Z2Zz6yGKLr/AAXbElaLaIfEltA/T0xalkBt3ljT7n9tn3XxqiUe27u
+gjLpMBkhz85mzbpffD1IWPRTTzcrouuGpunPs0VthGJwILZVyxH6lYArv5AV9YblNXbRi/y7++w
azBoe9mOVxhGes9q8IT6Qt69XpsisouoPgkVAbWO6cYz+M+KVfbzeVoicsfZhrAHtFyLdWu1SiyF
mn9NCwE5+ZGDq1/ndCl0j7skfb54z0myoUN25Vn5t0HqpPQPrCUK70fbAP2CdU61lo/BFtXAP4pr
LIx53sdxB0ME1VUpSyCDQBumrA+bfzAwXRkvu4K1nB/ydJz40Vmv99tNvztWGXX3tOoGyfdgx2El
L9bW9oGrVca/FLYx8H00VI8T6v3GSFThV7eyF8j3ah2mQ9m7icV9uyyUxgcNvm1I/Xna4mkr50iT
D8VNE4E2PjKsv0VHiEWi8l0eMcEdHsnKFFsCsfjH9hj/yrjGTpq8D5rzqwi4IyEdRZ5Q5oyTOv9q
4Y1TB06DFRsLsMI4ncnm5F0D9TGek2t9Xlw1ddzZnysfbL8QmrXdoAYi27SVvk8CJRFzbPg1sLVl
cIxK+ErHEiDEkzZYehfev9gdSyHnLtumtJPumWv25mXxokV0g0KHydJmZyBnNfdmPqpu6tYIR0Wc
ezR8uPh2i9UbHsC17gdWd7qXZ7gqnI0niPMM+tg6UvNE7K6Ng1yd6JDvWg5sGeO03gZCRaxLsClG
PeeiIIBo9waEHlQtvZUqOw9RMj8OtPk+b8ViiLKNhFNcE2x+P+xdjA6zoQl/MYko8cMSc5ExmEzU
hM4VYa/Fqm46KhV9R4oUveoVPeNkna2XhrFr0swj2CjE4MLOTFKa/DHr0+jaVG4kfAb8Ob2dNIGZ
0KbhYTJTPcneGp9SWcGhV/tddpoVhRJGEAl7e2/zjzsLf0J7036vjcrDu5BNg1vTFCwR/0HwcTPB
lSeCrBYvffh4O04f/PEiyz7WiVINxPuF1BijwlruLfjo08rX+UHKev7WApcdEF+X1mccsJWl6UyJ
HKGPFv+6xas9JAxmgj+bLSE7+KLNYaRU1Oxa4OLwy1VJsXb7ATVc4NQJkdojvZrzUkF0ThPqtcp8
Fioee1OagcmxLWvSSpsmGrSF3Y+I9f8+K9rKy8CeOSxsIriaLIi9XvjON2Q2p6j87z020/ljHspE
PlmrMoApfjAK6F7G46udDP8dEqA7sQhkcTAhtNPcjf/dwty0IfS7X1JeUiCgrQQqxO9grPJwkvaT
5RvXva5tJ68IHDm3NgGbRBhBTfaCFa7fz/b/ejz47kgJ6Dkm43QcBtnp+3PyIQhzs0sqLYc1L3mF
+Vw35ZAjwvpZxdsEwbZY/99dYri+G90GqLWl14Oe92u3Pc9ZM/66vcyFY0kSQmtlM0IEzHe0j5SR
rR9C9JXhacLxyZdj+jClYzKJsqD2b/tHMdLw3qeTzzQEoaVPzrl6bcTLTUC90N3FlWKTN6XiRjJM
kgdHdzXauLNv/7TdW1gzyjyyTaHxwcusNtSTXIH3kSPi5QFhGJeVVsLToi6ACkXmHCLcQo0vx8qH
hdbdzl6eVatEcqzHo99JxtKIVgAVKA0P9tnzsRc7bTnJ2HeTOkzuwWEAUq6T+xIWc3BDOKPQrrUj
JVr+UhKWY+fGLfjU2Fe39/4oOw/Fgf8cQ+LXzyS+NwaWthGxIeJ+O5LfuTW+PIILXI/cOhHtFp5O
VER4cLDP6whcS6IwtXfnQV+ZgH0MTg1MakmzPtpOOogqlc2WukJp5zkLRHGEi31RYoR9zme6NLry
GjzAfCgJFntFN7NK1S6e/mD2y8S3F0S0HDa1dYGHcBpYln/wfIQk3Acm24Rmn6diDiGXBZGe/S2N
Raw8F/6Oan4cCJXmHbJbyDjQuvlT4Vc1Enf+qoOLJIF6y1VPCFgBp0g6dvVjVlot1yOlNdwqfeta
U7ECnJMFiCW4m5/TdSXxGVQtZHlVaypGFA9qTSlvG7tr/hTeHtBB9zaNgzki4qXfBzwXZLLBYhbB
/8fa+B272/FljzYhqeJQEl0D5ZnJIIbc4OBl9U9s0g1BK0ZdeOfwZ6SgK+7oQH5o3H6JkT9OyXSv
RYTvBFzSex28QmLWc3Rx8ryAhoalLC9rONqUcejoHUg5Co/oU1FdySxYs8Eio+4F741/KY6bAnEp
LuGfq/PeyZpY1SuUWm+HIbScexRheqRs6WDDjN4AQa94YnoFhGZwTokBlp3GhSvmAnx5LFUi0nZF
CJxufoh2/DxNg2TAlCJa7/Z5nIjbo4ZxJ7kXKNPFvu2JJc4Tfc/K87EiPVsO0qXqacktMMLwNZPn
GGJEcLmVwyZsu2rRp7kZKfocvgQKzx3kKLo7Xzu+wGwGuFN0/ngyEpBeFQtHPndTOgG7G5CkZdSV
6kdo5RjUuSthnkXtOklGPIsCKcOxKi5iUZ7G+hMnvpFCbdBAnKsPxwG0afwAUOmxWqOe0PCzV/X1
aURFx6Hwi1CGNv4qH31t5yEe3Vw5hOrVVfFiotarlzxd1obZsUtVgpY+VSzneZV/F3zvyQsxmUVd
MF0jpWX8FyoOA7sGkmjq/JcYxkH7Kst7NLcvU+kwTdPio2mgKuEbsnrInTUvQK+SDuTfMNLJqswY
UMSEis6DhLnma1r6Ve0hVjHde+FxtTtC5Dxgx9u7XsMq5ClsUbGHuh99YRbLy/TEgPTzpM3v7eql
rALSxf8N9Xrl8DORFCLyyzb8hjC2+87oKsOzKMEgolFdfU480xubVvdqagOOYZNlcVUo3BKYunpJ
Kg/C3QPxwpCIS85taKar6BZUGUWmo5pKSimRNTCwdgYHYWU0ly03GzuzwFTbNfEpApx5SEMWZn4m
jXPk5oNri6nf6CAfuzSYiRfmL4hyrvYsAQ19kmtZJhkSFfDYzjycT92m3xqgDBTURUOVDQLlNsXQ
j3/DphCcr3URXUGVpI5kV8P06AE3CNtompo5apCiuPGLCq8t8s8+gG0AXHvPUMVgztevbnKX+0jC
WCNjeRQPcL9pSZXQEd2WXiTbLXD5gi/hF1MShN7Glx4/Soy1OsoHswGB/ezQQj2G8rMXpDD0nc19
wzddskhA8pWRIq+DJC4gYZwDvuiVE9K1TPiR+1FUlP+9wKcugwhLO3fJQ6k45vgHP0Q/k3pNpl+d
vkrAvy631GSTC2rMIQ8CKC4lPOynnH0cmBDkX7XAPZX6tDBTsYr69VqPKxO9W/7+bb0B6hb2ptbA
QBRFjRLje34AQdLvAcQrL7fou0XX3nufu+O9zXGO2esMn/mAnx+B1TPZ0oiHUQoQl9xp/eEF6pCm
OpSbV4rXgAcmhk+AJR/U6uYm+UNYn/M5tuz2y/tr0M9w/warRU/x/OW/R4X4JOiUlTM+3TmNPTUR
H2KQQwYM78j5KetuAWTcMxd19Ka87bqUdn3fKFBN0C0sV+tjcUs9Ys6h7/IxgjFLeJmwwrLxK3+C
8HlQzUwHG5oR9xKqHaXGweFDvuEsnXKK0fbu2Fp20PLdUFXsLnArg2F7YD13mIU7Su54KvGCPLdX
yzleH8p+O57B8PEVG8UsnZvr/g/JP7vqCfm+yWsfGBSSlTLuiN3TsUAh/sRaYUw9wUEVmKpgjwdn
1FS2FUp0EpFHiuW6BwgNazL8VrxNpkypd7PWdd+eAlhkMvmGyCH9Ojf7HpLxRw28GASkofT9cXtq
kJRwA+mwzW3EpRx5LhMQAsZGuzdSIpwnvAvbmxyfu6hLIbpPHmVMNw79sKqze8phoenHFFqeqacH
DuI6FZXI/RuCeUmPid/7hiqCXnTIcV0jiRMOAsKd+TnfsZNlaj0SZOJEZmDcQiItoqW3rmSISl3o
3CXy+WHoLoP9WkmeMhSy2QVrAQ8XmgwjtVOzV5CEJleX0oZISqP6zmtbEuOpT3yEKJtARQw+xnhr
mVCb2VtnbGzQfaf7c757UQHQZp61oIkq6yR0dmGXF7ufZVAY7eXYu577GOB204YbEIyELTp42iop
qPlc27dUgx8WnhBcEGTXyDUJGr2ioZ8Tkvu+xQCbpeREIJg3m5Kao/DbTSARiWSFn4CH8O04TNAq
muGbTf0/DNM45ecagyY33xl93hLcdsgPvex1xVbuqFiwf09zAoxUYlP/+fhEgkZUFZY3m6fTrb0o
WzGiANDc1Sqe+4uFM+iXt7VPor4CP2cxoU1jD1xDuZPhJYQaBvzSN3xXivzW8K7Igzq0itRADpVS
IWW9KemcCNE022t0BcpI8/9EYktTpaVjCXemmBxVHbjXs5vdy/KKINvyysqIXIhMEqs6hudT1bJL
dii8r88FQO9B4lNTLdL5wiUTcz6X6ZiqTcdaiKktJSXJrLbdFYMWWAgdyQu6yV3t6a4cY8pME1nJ
f62Y6duqkGv6Kn57vf3xHgsTYfrVqrA0I8M4XD+476QQf8hMAsnTADY4Cer5w3f6bKz5k+QhtJ75
lYukVvExLLXkdJXxMjTYJC8usHeECVLYg82Tg7S5WpmOJemKx3ySTQlafFEHwmjbVVscAEGztlws
qp4ClvQKIDSTSRLnb/F8XPQNaLwLz/1FfgxFKaP0jvvSOFxskWbLlmo4Laf0Ak7IbIMb6/kPmSE2
7oDRzSrw6qAuuWcV3tw1DM98N2jGVKLDqfapfK+to8jSY9svXLCMdokPUZyEPRY0lJ3qmxeWRJaL
DLZPNaRez/F18Dt0q45HGRbepALVqQGCy/yr3jhzVmSOdqU/ZbfiVcng4WMoQ0IHmzmEG5NzvR3U
tQKR8qR7GmG9F77TwuIGMOuoCb96/MKXrizvW/KwT9dHkPClYoRrwreL9LaG9dBbCxOKaMym135G
rM/iLINOQgzuaHiwMuKywrb8UPBkJ2Rvw677+N9P3p6TZX5PxttFdKv3bNHKVUfDIuzVDfmyCco+
ZThpgJGWtAkG0aI8rYxD01w/a9NFVIsiLmHXQvwjFUmgp6zcuOJPY4Uer6Ska3chktuzPqLbWjSc
6NF4ISkGKG94YerG8mhGr592FTw6V2IRYP8Fci7rYhqTZNL8CO27c5EB3/BxZZxpmm8VmZPPky3/
jc+vStlRBLvcD3eufdplJcrxDpDCSb9B6w5pnoMWpd09qT+2rZf4ugFGCQ6RLZy9PISeyCdB1Wd8
A+3LUKZ+Nh8TpboE8T25aRc38NvyZ0v6/9MbUqcgUPr/EepwalBpyezY3ZsEi8+gXxO4rRBe4yWw
G0cE5FZIkPBE5u9ZQ4MuF6ED5EjFhfURg/JvA29DM+fnsXGZeDF8BHRwSrQZZAUgO9cDVS7rSC1H
Ftk4MMcInPL2ctFg+nscSQnmWpcZDkZC83B9bT77MG5TqwQ2UZbp9OtS50cP1gHl9flmasoOsY3G
l9ljwrCiswJ8tMxJH3CcSMplh7ebg34Xx6f+ieIpt+UZI+XKoadzRThkUnIoaoGz5knSfXYgck2O
VXM+AiENQQNBVPKx3ZtMu5vwIMDNXQskvpucaX3y6GUBz4ljuWQ5yCL26vPn1y7G3tHdh1hEkKd2
elCM0pnkTZn75nL1/mPzeVBDVNdmtjSoq4gbcvRhboweBZmYFqIrFAP1f/MKpYgK6+Ul2WH4hfoa
MH+4BFAmNr/JAUYjTviZuxSqKRtm5QzYUhJWidiJwjnKEpaVuFg8QwE8Hiv9t0OBZYla+t9tGrPd
RN+dj56wdkqpFaOdnka4sZbiRkBszXQ9HONUw6xmoSueX3/YxEeUxa5UC3uz6gKB2IRVNit/aPO7
qaSalCqwwrbmc/+NcIWAvRuuIMY4nUL5QMXU2cbkLGCQBcRTNWSDOGDivnMW1rSkazCiok92G/bD
2qbA6LFjKnBgsUHzfHHa/pb7gT5i+Xtn+QlEnaGBHq5UDFNE2yujJJGtJ6UQ89kXRodn9j3sLX4z
nFvt5FnIKQKdW5XVSEGsiSY1qkkDZq+EqUD6hYBvL5U45TYlZVHtVuacRZm1/sSQQM7XBEYnWYA3
+bFnZx1PtGMlLuOceNTmvAG9b2DvO6uEQ7+jFUrXxk2ymC3jIpZJS2arNEhWThQmuQXpjDi3sb6F
k9/zbeHw25LMhpr6grKoP4o4mFtyroMtLddyrohPIm41I1oLkoTp3vrIZspdjeFwWJzybNd1UAjo
I/PkIQMkmmqAOJj3vEmJNu9r+vz2uInA87ovDRK6AjLi7Pqu18bHFWsdSu6p3bvcntdj4MB9Ql5B
HWedSJfrNvSTn0KYteHP7RI9Na9qD885tVyVZ9QvB5taFStsWSRGDfZZofcmfUaAEIhjtV8bCzpV
c5B4hXR+U9wxPZT3H1IOnjtvOq82wEV4X0Q9JMe6aKd0zGBaHN0601govxfL0rBF582Vb0Wysf7Y
W7GlyK25hw8Ycx3AIRPGUP6hCFx6nWjLEmxO8rEfxwcpVKGAQqDdjvsrstG/LAgM5qxOm8joSwJP
khNdnIb7s4mzE84Wv9RFTRYyz3dHSxnNdVnUFE97NQLc37bLzT5Hm6idya4ez55t9kc934BlcF3x
hEPonTalfF01FpU3yD8q3awYWweGRpux+9XOeF1UwtPp0NHWq1/r7Uyuw8uKuxzcDHC5Xv/IvDEf
YJIS0W/Sz9l8pLkn5z9gmogaOXd+sY611n3zjoqLC2LLkk1qd73o/rdlJjKRAyk3iJSTMyUuEYEQ
HDvJKLVh4FjpI6CUpg0Se3GmRDXfRDWoDfgJ8RRM41UzoPQrrLwJpGKoulZukqgyYm6vwabhyNYL
MGtGPlvrutT5U6jHMDTnefelRrPT/QX7tKOQFgpYwU49lxhMX51uDcfItoGgwI4R60kCpPaRJRaB
rBDBkWqHhxBlSErjJ+7gIQhsUQMR+VpcrMpqbhuFUE8XpMJnItTp9cn7rx1E/PQEfL8UYMUA5Q1M
iR3bMgnXj4RqSsPVd6RRmbI5vLp0RYYbzJbNKMZB4oCSTdffEd1ksUq5piloye/nwf7lvXTsjYML
JthNZEZcbvgUdhxaFz4Ka3fB9lC22i/Pw+ns+gP9m/3W+rfVAab8klxozbOqnZmSrmqobHDcwed2
K/gSexrnqSxi7dS+uWxUDOOXvKEQwHYOemDf5bNMy23IgHpnqjMEAeEm57Be5Mu2oUBEu86mrTv5
S6xKsWdhv5JmRe9fDhCPysGREwKmZ0Nj0DXyXb07EsA/dApZOtuQzwMZXQfOXiA8mTpeXBrlUYMu
0QKvvIVBLcAY7lu5Q7DhSf47lgB15hVqcHgcfkZkPAe0QBixu43l6eocJTFVnZy7VVVrymLXZvG9
XndQGCtEVUJfscdR8J4LgnZUnUOUBkFRt+4gI0zvbxYg6/xHRpqFzxBXhLwzVmVAxSVGyTX2T1/j
XFzrJBI6EucT7heP8RefqfPnkIEcOAmbAtxy0CXxfRW2hbQxOgkyHW3p0OtMcZ+F8ROhpT6UQhUh
rFyA9fSXh+B93rLE0rK/QjyeVg7MgLy3/6NAfcVuiLUyQexjQbpwGtHJ4eOVSRQqaTbbZdO+M4sV
0DvFDuUe+8/XJ5KO1y/p+3tXvEMQxJnj28STkW2IwrPGpk7z5z/ib0zYicIRsA7WALNJASWPCm1W
qcQ3ffIB21LS+45vn+tGbPxkdEIr/ozhyuDe9Y6ZWopxtVpWhyADW4Z/98MMXLHX6Z0lUyZh6VD5
ESjMi+tgrEQMwGP5jKm4XMhjBtXKydC9wNVKPHGuIilO560TgkaU5JCfVUlICA+lxRYjQyp7EStv
QPmmX6EwWqEK7mcKrzuUWSepn44RclzeSBVeF8VLxdkmqM3za4Tc6dmBetoNwOg6SLMadGswudGm
in6B5BqLGOrmQhusMBQ9zHjYMPH9dyPF81iA7XT/5/UoB5TmttxxPow30/Nenga0vxmrIDTMSgfH
0Ws96ZRYKnHGb4Si/k60osDeBpShh78CGuUys+/w8Eg89QK/2ILJAoPOmDtWpHUk4B9DVa3oop3r
dvlK2f7p9GWpNyPv3dVatKh9WxnAaPS8jHOXvcD6fJVMRjXn51rfohxy+WLCX8ycAI2skq+EgFpI
ryY7RxsT7xEFv1edpi38iwpaW4uVbXcca8bF4IGDUZiZlNVFzcpFdZY7X/H0sALMF+yq1P7VevjZ
jMqBNfKgG2NX/LJedejx04F5PCDRaGeZfqdPZqGR+C26SeyK8zn87OGewrtXuyarSnuHqRYtFSkM
u/BLSWeBWAakAl7GypuIVTB7ibqyrbw0SLMf5xWPlu8p6bs657lmsYMHH5mEL2PP5i4aePDKGhNV
PDGphAgqJh8XSAPrNZ+JsYVUGrZVtTySLd77DTPvF7aj10NW5QjrEFvIMbcX3tAZo+nS+ydK/knh
Fv+VJmR+tLq7whK1/aP7I31BAAEVduUwa/IiKnxo5qWadpt5OKL7Yiiu18rH6wb6DyqUP06XCIQB
iYv0+41WBtqm2yRLqdtQNfFkX4nHFFfjz2+37rBsRCxRN5Kc6lPM2PWtUu8KBXp8dLWnxH5osTvJ
sS0rJLaESWvIz07ifPSATcB+Oy0NgGINKg+HzHH73qGB+bn8wO0/w62W9UWjmsg6WwzacIDtgqdF
MguQF7iKg83H9HRw8HVXN7n1Jgt5TPLV0ushlmN9B4SzJZvL6f6W61URxGPEHZg9rNPSKwHM4EJf
F7n+50ShGBBeF37zS0vHhgw8aqO66E8ZENQ30iWDdbjU4//UZg+Rj4BUUYMo9fjMLGb48CgSXGC+
P3+E+VwlE5aGzmm1Z4djzns5FnlUZcPVK36zKo5UeXlcrCwsMVPuSJYzu7rmJKvEQNtMqEM/yq8Q
KqMEiVMg8CouLF8rzOxZVFTRFRgY9kdM6zLQEp7PXfPRi/F8mzC3Dg+ATj/GXeP9AeJJsapCYsow
/x6H6k/wgzEau7QSNq80X2MNaBS7RJ7q5MIiorf200J9ONsswuBO+IdWKZZRFImx1xSP+QuOQrRC
fGvOIDnhpDv80pXOwsjfIo3rXLfn9dJa/ePYe4lz6p/P/1IOcK/oiRX878Zn4r3oQwuImJQ+YjS4
u5VqVAa3gVOdHC2x4XhV+SZR7FWQBZeo/NqqGIf7EONDUWXvrB87PdYy5ptA1xsy63bPkbO2EKry
Hd9T2a7vQgqf5VPOntNeuYSNgPGrKx0hlnPnOsLgucG7VzJcg3Rb6aYOLP9b53JlzDads3uo0B+F
Mc+Uc8sLS/iWKdg9OjBukbBs3HaDzfe2+08+IznVWZnhM4/PR+UQoEzxhO57FYLW3Ix2bnMmGNuG
izGiirelsGYth5eizH2/vn/akSd5Js8GM1Cy8nGMlIlVPeHwq0CfS6YiEh1qhYn5iA8pJ7MVAlmS
vwzfaQaORVwnUiKqSseFq5h4+UtCDVfL8ylBq9L3nbKo6JsrJTE2jTafhD+PXrsmB6ymyTgL3oqC
Y+lRJ7W5SPmYEovx8XNkbwr79D65uMZK3v76ucxBWwVGGMjiLCil9XaBuy8a/uyuZ3POvV6/D1Fr
OY7pMO1jtpvEEFWwbbf8x2ALyIbmoKkqzi5IPzkpUeEjtaNtMZbpnzfQKNHtjtMSWqFMxsT9ylLA
pm8GyZvszAxnjv+xLY8FTzYcrR5eYNtKOuqRtqlp8QDVvf8VL8eSkz/NawbZooLP6JiYO6owWpJr
nmdTHE796epvPAZn+dfBTIVBFkOJeJEFyejSOWti9htUuYUvoJQLb0aP3c6YzSaapK4Kv69FE0Ip
adt157Lr7b0/AojaJ2xqFXXqIEG9FIqzLX5yugQUFCFqLypPpl8eiNF2F1NbsySv3DSNo30gEbDw
xfSSgxPtLk9KLXzHwwbAc3vAOO/f7bjSXv5Vx4ySS4qf4mToRFvAAwnOQsuzIYrznd+oNtL3P2QT
dxj+YLhuk/oMDl27vjQvZNLGCdKzN7VxhsmiX6RfC1vw5JdF57yiW3MVbQ/KCaT0soc+XWRWEu3k
EQiG6GP9RfLvk+gXYOinVwx+SjtM3Yc49teLRQig3qhpceIk2nZk9IH4kYltyzZRAAElpKKBZBcI
c82YplYUbeTVnhNJzF0JhFVyKMftzKunDnUVqVYAr554lyBKVo1ttjzEh+jwMKW6IEL6IVBa5g6T
eJvi+Nl548XF7ogG/gEMjQ6JI0NHzv6XYNWTF4UjKhNNG0I/yCfAYrGyw2YeGqbPpCMB0TSJdnZD
YzyYpbp8Lxx+2QbTRF4jRD0pei/xYAi4MpRyuBS0BusDATEiQMqheZxf2as5irp38E4pj1FX/N0u
H804dd1qrc+bTVinPMkAJuPCEiKUCohq+bpvA4ar7gjQbIDSn9jYGjlgEnv9gCrBlimsrY9M/38q
R7NAcAWK6ZXekG9aoHg0Upk+fud3E32EipuWfdb2+dwxKkeGmqNu0pWjkrbG1G/21nrfZmY45WXP
n/esBLnNivxpgFwXKHWAsIeYF70p3SOC2i9cmMfM8LJNoWa6+Rn1ooDJg6wVAxbUEazK/qtM4VXB
IYCGWXADJYpLu+ZXmUgK8k8Nh0t8SFzDAL2Jti+fKQuAxYhSkpoCFoEtekV3oTHI6N5jYHCEkOKa
OgIplsPDr2NXBf4Udal1Z+cQIJzDTBUJQeeEjQN8ksqLFwWj2Q10t1uH1aCdLf6fLnUHiRpE7LwG
o4QxFtJeeZZQoGlsuCbgPJYUtirycJcEbDYKfFvWpsUBQsEzh02QAcvG08iTmPO9hW/jCO/9Qx3g
MofdATW4BN+zb4qkU0+erKFi1xAjKE3CGOEpLpzAgxq5uTm0Cu/5CT2Ufo28IR08QKc2foy/CWQ3
MdixtpX0WcIzDF92EbF2FG2FmKWUbiC2n28zm2TN5x7TI9i/eNjVjGzEfV1M7vKaMZovfqJRgLKH
6Y9LQnsGrJTHyqENoIZeR3/dRPQdMIw1UuizI4t0J45MW8bxTCt6nUK1T+RJhLkZNZclDS10hp9S
Wl69QjbWHTdHBesnwuWmGBhref2o3X45uF/RoWO/sP6/9x/N3BHIyx1PjufBtdonQmnsDmzQheFV
EL99n6/Fexbn24OU37EEVsrJXNjviB2B1RLQF8LcaOHm4mfs+UE2na1ewjF4PmoxFAl8XqZHwWez
LjjuKajFwZVhbLD4v8VokclT2jYPY0YyySAXhOuqb3tl89XIvMB1GlQpgkwIexx2bH+AUCvBYeAJ
bAZ7ws13paaBnGsMbK3P9N+JqTn5QEundm1dDnNnSxH4VIu/Y4CdfbgtDhRzuiA6kAdNIfpSI2Op
R4ShlUXIjss3F4dOvNHF1ZuH6SHWrmS2ZLHlBo/OwzcvTuns8H4ijINbqtDzkx9UTBcSgo0msvYO
iGZRCt3IXI+P7Z6vQld16VZkpFPQlCAec7QBxO1oIwmpwuY4rAwQK98woeaEa9ua2wFXTbw/kREs
xi0RXTycx+GV7VxJ3Hk+MEubxScZ582R33b1t7Mfnht/yL15Czk4Wc97DcXaDIXFtb5u50e2wEk6
ftWMxQHhWFgefssG0XO6RwHQ5EWkx1kSuUYDiGFMA86TJLbTYkgTvJsRRL/CdO6Ce41jIt71e5Ou
3Sr0aWb9NVsy1N/XM55EM4K0g86zGh8legBHSJIy4QHCgf0ZliU8qeEbMa3BTpusY0ta+QSwstzp
kg0H80bG4/RMZp87y9YDel2bDC+bog+zSOmSGeiLCFBH+oafsd0lIaAsrQ4pChSsph9bXGNCaeky
FEdZe6YXae8KNQx6zDVcOZdPyrnhfZNT8hEVNrlr9rh7iSa7sC6QqVpUZ4Dwg3XiIyP5JYij9FaM
/4DCa/aKf5R4Etxanp3h/nrV7dvJEp/RvbM50vHAl/QjBea58S2GEZOZYga0Q4TM8Sk9ApZfpxXM
VoDTYEUp8PUWxNvoZbF0UaPQynuvyQZaYFlMaMaWYZtRHsm4SXdX7yc5GW9s8+CJPRmZS2Xc6kFE
3sVqI41mZNKuSeXY4Huq9pgoztvERC7JXTExfHMX5z/MBPCjJf/xjYj40lg/5yPQrESkdo7Xfeno
Jj6KdqYlQWu196fKOgmZ4tGzcNTtYPlZ+oKslY7pa5imiqOlFjKpDPoV3pQhKZdXp1eRCgWx0T64
bXfTmyJ8wmYKW07o47l7qPLRLq9R7zIh+YEr0576b1yg1xnmUY2LGvZZJXjjumzC5V6GeR9k8RxR
MapzTovyDdwT44Edma9owbQoTGORbSW2FamIB/5JC1xRZPEiyfhBBKSco2UI6D0MA8V8YHjFO3C2
wUbXDo22rS+bfdEKq0YU5AAUWW1mUeAqpzu+im51jAdX/jID9tdH1TY5uzSQpQfTBka7rWeExE+n
B+BzS6MS2qRBh2ts6CViUOHRjgCqxn5BQPaGip+TMR9Cp2BmYmFCW7GlKJNe4NkNdfgo5yCrrinB
zbwALq/x/Akwa5U1Ogbo3Gn7WagbRqEvdmjLg/uC3a0xYmh6dqRcKKVke7wgqsg68pY1+FFUy5kx
91b1XnSSaRDHY1Sh2lvc1acbkCUv8Fbg4upy/oiyX/70O/WmNdiA87gHlivzqPPM3yC/S7pTLoeT
s2hLp+q31t3bgauBJk1DiQn4uAUOh8bCO1AhUafwdls5GYsAZMLKcdVKd9RSaocE3LJsSByqu1g/
m6QPjjsO2nlJsSxmGx4rlHxGT6mNtC0oTq/s/X4g+UFR6+Sm+yicR+XtZed1PM3HzT67h4Ag/epj
oZPTTwulpkg3sUR90EXk2YHHl/xQ7UI30IrLiuvLTXFt0p4dLABkAuGrcMadytcU0taJVp1Db6ae
MnrzoDnvKqaepzJJfY/rIGgw+t07lmHMU898OKNxd8pgODYL//3yWm0KDiRnmeK9LWQki1OhxD24
1EX9Lgzg6LBoYqAHF/a+eyHg5SuJS9A3K4GcWMrQuMnQWzjlPd+1pov9KyV+flkdb+3dnNYA9i2D
TD3yAYHcx6qMyR4d2nnmvjm/lvW/ba9JNE6Zah/AR4QHmhlb3/AV4iZKfVj7rszL6MyiUbrY7pnH
O9h5AL0pbjDat/H0wo3TVyVbSr28EeGQEYAkwjJx9vM+Gegq73MjJoltZO0H5s21UrDHbJ0CEgbs
NsskYL0iu9Frm+PaPInc3mMOvgJ2VXc7nPDKK785PMAw41j+H4ChGoBz/e5omxXzc9WcYYjbvYaz
B7UBJr1z1uXODC8NftizC55lQJQG11iuFtSATyN1mNsRh/cTUpOCnMWW1k2QpomIgwKl/4JZwajx
fPY72FgQgRgy1tOe0yKilB4hUv22M+8eiT/uTWG60dlqgYpG0svo8PTKK3Dv1dAAutHCiXzOo2YB
V/ZkWc8/0taxgzHTJ7Ws49z81uAfEWK1/UkbY9EDSfpoRn+g2MlOsuMN8oPrZMLa1q9ns2XPKl6x
r7kkLkkoPBKvIEg0E8jbHHmUd83eews0M+C8JCHGV2rL7/Zuyk4PfXu84cds+P18JBl705bHx33w
nYr5zfzXLLasbQ4k9brp2QKCm1Kzhmv1SycVn+/lRLAu0EqTd7yImIiMb+gLCTPuJqixEOmyvgVn
THQLYkVcQ21RRXebyT0TfShBEcNy82YI0lgCI2fJeuI11KENrphnYWoJ3GSEXZlWlrNhkcPZlp/a
TCQVaY0OTM73MJK2vW+4OwJkb5HR9yP80b0wCGsx6DNalQFEl0DheK3RgUlcG+LDNr0Oth7tMhfe
OI+RLbzDAhsjwOXJhRnFdfoFhx74C0vsWoe6iUOG+XCd59ZPILQPnMX6cPGaRwFgg/rsgqszuZLY
AlkytePyXoKPXePK1w6VlnWqqXxWLJQMS5EK3/g2OgTvHmySaHSdlmUR6pdcA7N/cycfB4kEdoPI
OW7WtRYnh12jebZ/zFg+xaDu22zbpH8BSFSqltL3E180fOKK48lIDrppflGdxMvhilRYJkHj7tTK
ZgRWSpTikF7EtlOh8m1QWgfhV0FQAn6RbvA6oYdXG4LR0TJbaJhOn7s/7aj9IIjirnupxd7twrVr
TyYxYvk1mqDTIo7BMhmtr6jzJWWb2wiPib3K73EvplG62lWjoYKjtcwXSi6FK5MaNCdApCRRUan/
KDW8dyrU2pZG3YQpxl31LwAZKF3AjVQaRinjkF/foUxxq4w2LUdHRg8DidZz1uP3btj8QGlGHIDH
YPsyz3vyUHcg7Pq1OSqebQCPgwIrSu3mPYOAUwAo7zl6DEuVQ7ctO8vBFOU8DgrjkKzE5W7LhTQy
sW4na/Z8qecAVw/sGWgaL4P1ZieVkwXTXpW8TxcJXx2wop6UYCYG2KcnYbrGPXavcc/VVpLnpNnc
GmEUnQLjztuFQdNtybfo5MNWz4/CDrEPvDkJNimj9ilD1LhcxhxUzneMOznTCzY54yXvOViEeIhW
Va6+GuX2Emi1qx9rx5dST9M3nmlhJ4cvTHF6Lo07iakZx9gA4LLMzL/0W1w77hilN9yxn8+DbqcH
m36S0zTedvNLR0h5FAd9ZPviDWI7qUxC3yEx+9eYknQh5vg67ywCXhulcN5DgoBLTfU0N61+zRq0
ERT6W0wlDFEvehoMMp5drKAMvq+WWV/MY0QgdW/e3po75TILvH2vwW/utxx0zW86oTT243Y3n0c0
qdcv6a5T2FWGvwTVV7QrnOrz+9UXxbyy
`protect end_protected
