`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kon8OECIONKeoKqT81Fz0Gn6vbI1XpLQMw6WdjBkolly3OSseR/mfgnhKE5+FhP1oSh/v91OAhtg
SVCnw501pw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d0pjamPtoTce3pVFWeMgtstHxxEXoxZ1Vh6p1QW12nf6+/u6bywAHpQjsdyFpBnzlHgja3Jaufbs
nRwtGRC4MYso2GwbzSiMq3FL5sEHHfMqpW6MU2LC/DEhpEcEHJizS6Mrx+qje/BtJptcCNnzbawM
Q6RWkjJ+nCKBD3aompU=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gW9fqbfufPNBemrHiMDyuTTXLE0spHCYj3aAIZyaqmsoDxm+pRhdI9tjdwSc37mXgqNHdaDXcj3h
2JPkkHywbQIE5Qpx/gro26hrYiV8Heyq/JJ0803283ZtLc7PaS8KMI6IMQT4tAy5pl7jVjHSSFWp
oYenVVtTY6tOqaBds9k=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ffQ/JEFlFfAtDO0OHjuYiGGfe9cSP3DQegnPoFmdd82eO+YRMqyeNGHBDH5ZEON+W/VvUJDm3ONA
Tkwi84d27QpVaWd9YiGp58sMon4klLW3x34n1fmVkQfZzSURo5NhZCiPLiwncl0TQ+XLtzcWxr8G
gHSAIuo4osV9bnO2zqjszIOlZbo71v8ZzppGv/ob2oszHhIpUV93P86tFbZxhgaIZ5ggOc3n6wj7
+YYUoH0qooir0jnjAT9MZbgOLrcJb7hj5dNNATGwZX+GoS2482kMOSs3HTIyMlPEJd6cK/L+WE4H
BedJuaTvUEe3plJ80yNZv8vtkeRH7hDDIVp9YQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RkKtRQT6SauA+4Iu72h8PcS8FHstLYHtMQv8jZ8qlYfQl0p88u7HV3oUV+ocLUykJbYbO0dAfidA
tl0cNgdD7wCki3q0aXGecZifyC0Fx7IFfnLNVafC+yKTpy22Mt2ZGn4IMyEYV8Vo+u3BW+vN1iWN
jA1mzYue/nw5gdLLbMgqHB/uyMcRCv8a9NmIzy1XH8Fzv/23IY6RCGIe+mu6wwzfJz3GTsbITHUL
O08ugqWUwFG5Ara4Ejp8h9iF9N+eXX9MUVVhTfxSVfzJAQgDK0567i88Nafp71pdghSCJujSn/yX
cpZtbl6b9wnSbmUmfEDxhCx+D38/REUD21JFqg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WPkGRJB3diVeEkigCgmW0DAqMnpqZF0dm5AEsDTjjqfCWvRg2IrxHNc40wr+nK8rTr+eSZ1tTON+
PA8k1OWpi35SJQ8qXsEOVFLgkWG1JrU2H+FdbF+mJwm1D46A8op1LazhElZ3io1oOw1Tnhpsl8em
vME2tPnp8vAsVCrLwMnVhYW2OnV4uh4XykavqnFr2gFuPdnxaF5SnHNXDOXdV//9HuImYs/HOoZ/
Z9G4BWgFS23NL+sURmsBscgWcxaxsdjYL1JpkMx9trjf58YT9zJ1FWM2emt9TjmYupggjCwRYE4v
hYr9LgAJkYORb3SI4msPYk+U70x67OOeBJMwqw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 67920)
`protect data_block
3FivVYWi212fUIjxtQZaRql1vUaG34NvZXzMevTH+Xjn2hqL96OPWWB4iAb+GMvbM9thzhZHbW/Y
VVspkeXUgYgWxjfDkIlY8HfHbfZdi6cWlcUCViJZ3gffZJUgM9lDR5dnQZq/ZHWFimZyqBGzBVcf
pQKokNFnuSRhMZgctKPC1PJh0BfM9HNDRCQHggeSAR8aGYw5NDg5onM65sBcOEMs2WThrJzF+be0
oXZVbBgkFomXZ6WR5YX/9vJRYDFuqJHEQNrUImAKcTT+CWws+BWNeHDyrntea9Dof/OdEhAqX0Q0
CUSU/fPujOeohgc29bA6qIbWu3AQ2L6deUoq+3wMYJs+HSIvpqq66VVOVZLcU3h8gR98p4RARduj
5MFbG1G4rlVdBL0lE1pO/n15W4RSQ4xw9tAhQGDEA+sTMGU9LlG30xax5UD767KeMDgxbxKRWV0X
4msgnEAZKkl9laFSjv66l52LlWO/Mi9DDr+E+tAQzIlfPZJQL+A0egTL/81x0/4IB8To2IfUHHNA
wxCdkOkokm43f9J9kq8dcmnzi/Kuj3y6Wepf5qHWTiUFmRwVJDL6Z4ajxGctvLbRfCwUqNCfjfv3
czlizkmiCalW0mILFQHsU/Ts0Dm1/n4lb4QW5c7YCM9Lbhz2HZUjQSNql4X81/hzcdD11Ibk2A1o
9KNEeRjUlIAKR9cRRMy6gxZr+UU30IFIjNIszxSBpFGXW2F6jyaljVegYmDgMwVTJSY5B6NXKnyc
tnhUTmk+Qct+7heW0R1eXHBSD9Ws2xuUBu0qFxv8LgEfpkUfr73BhLmDxioXVIA32Pwi7ZCJP521
XBIF+DwB/ln5MFG1sWuQnSjB8PHME81BlB1ZcRlGesAeTvSg5kjg4J7JnJU/+h0z5nfN5IhK1hKT
MVdCSdBOywa3J3TpYIEf7bePARIlFd7Q4MYR0lL8GzaHN1M+DOnUHGnuorAKThr4to9UTbtzSRsZ
ZrnmSRtYFGI2ivesIgEvse9Vcb1ZBxtZH1arGzPd9UOeA5mngOzlmL39pAjPdOIl7DSgbA9ZG6ew
qHJUlSzVM7AvAeBuo/cbSXp+ggma82Md0pz3nguDSn0RxyxBuE0C9jbDFNzAHsOUOPXdei9fhNTG
Ichb8bQKyvbM6LM7Y4/al6jY8MgeDQhyuTIs/boaLdZfmwGoGvj1Sz6+FI3XlKiR5b9330nivURH
krWxzLlB2ZiFoYGXhFad4UHTmr5VaxbC7nFMitqIZj4jsoeQenyu+6tUdGnhjcfSaAiOzkG7xDEg
KxgLSP+KjFGuJobm/IwICuEBXnhwzBmz9YZseA4PNpn98vHi4ooOW1PzRKrlVgRtd76Nv5hHAFsZ
G29JjzXcEpRK62hUIdPUI+jmOZYPEbhryatUY+3GyAF/oMRjRMig2Mr4K5kVFB+FwgxFDcOlq5sJ
KHJh92qdOJXV+2yDO645P7EtVS5tF8jdLJj6v0ZrNdVrWmU4AfrWwR2JLF6jYD93z+hhXgmGD2n4
uJ4oSho8nOna0kqyDIa6PE+UlaQjLqrDhxXFoB9b+EJmjdCuSPSpZbOUC3S3vHZDE9W2QHp1om3T
xxilSKF6YVuWbAlvnXZt2yXA6nH68rhWcXFPbLArVf5JNb0GGlhoHnGKK2jnquAsJ/o1B2q3Sy8U
uXRiHOv8Sr/jn+Zx7Q3fhAtcqQK0efyg7pzcQULXhreH0W0Bijz+5tggMeRdZVqmpTK0Eg/bZwW7
HyQTgJAQVlzqCueMhKgQctWIHu3ZrORo6vaojgWDQ9F35LooLE+lAlhncxDjDpebKrPdvXCdgc3h
AnC+NzbJKl5Cg32gy4M6hWHarD4PgNoG0MpipDpEWxrvxQQc73ZUjGflEPoFtMHzFycIF3UTVoie
iMB77oERb51/MzXy0Tk8q7bMsVoWCgkAfNPVjVNBA3NNsADq+CaBdIEOod1qbB8Kq37LXuv2dfJi
gz5XNqgFPuC3QXNaZsQa7cNeCqy5cixx3cVmfCHBK400rRNrOokVHxcGhoI6Fz+giRPUX/mGhPWu
8R53z6MwW8sDiod9Fmzasrt+al5emvyZ7nzwMRVvGutczf1RmmrgKb6nRIdAC03UBPqU9Xq3NyF2
CSjO12rVk92cEbXVUdT2Ja3geQe/3p4quzK6qEixtrsdjX8FhirByxCHrjk+GCaG6L2I5A6N3Tp/
8Sf7cd5qN4sGUc01JyrQMayLx4hisKBp8m9+0woVLPfa8r3pOqWtEY67JQxNgUzPrjvL1IJZ+xeA
B1aESFyiGcnCUJ3ZujymN9e7r1jJfXQfWeRZ+Gfazfdy2aO6utXY2MMIqEhUtPgld3R6EKm6/ub/
+Fhpvx5LM0zBwWNUq0kYno6QCxeq5lmRL/oHD8rFS08zeXCKy61i4Wy0qV7sVM0vP0SsToDYj7mn
++WwHGzRJJGUyaMYZWhtKuMF1Fbm+zMZPdCLlIXRo5/wVfDa4RVo/zXR6SXfyqWFRgPM0OtYww/F
pyoD4SDjZrHfBgFCY2D+AdplEIQdN5wacTIAne8yhLTMoOtjZ0G1naxntYzrAccYw4B8P1K/DLdM
I15a2x01tnaQiLVNbII1EZXemwrLvz5YGTaqiWFjNg0nDYSAOzHC3VpuzjgSHbWaQqDs7s4aOebA
YYDbzaW7Fl2Oud3K5xEtoFlxaB3s6LGRVskgTpJVTGP2DPz23/k1i0gn9w8Ndxagz1Pct/H7bspO
DiZL5abmVlq7bzhyskIYvMfzYWlwVrD+Gc7AMtigXvzIHNpZhsiKE+eTKXmOvc5myhB8TTLsY98u
5nUz3elH2AbaDMQAEGKEs2rn9dTd3MM06gWXymErlrUaRXoc4E+GBhrFQrAhAvZj1nGU3PxNtYLu
9wR5VY51shIpjhOvmTyAN3clBcP3qcS8FCrs0yEigtw4/FlgTa/Q+vJu8pes6j2qA4+DTuoVau3Y
0AZePDRY8BJxdT5sQv8Bezvj01fpWfVYmpMtKRoVVWmEI/SRMbJft+NTxeRKRN8TdyQc+C1seFBJ
o/dzJBck6CEhIyr5yWU1OmjgmuCuM+UYyJDVQH5bCT5B+V1J3pNn5P5xCNWvKCTm/TngPzLnSaaY
AqGz6cKNvhk+cSYLrbAruoicxCWBsS2V0lbVWEAN5rGuWX7NrIHffZ4d12EZHnXumqQOX7Ocm1fn
jK0YGzasMv3NJbKR66DnA3QLmhjsr2EHbqWyLQIhnPKUr5qp9BlP6BmoKy5NELrk/L4Mz7KNDff7
tE9gKfOK+FjFdBuoSSIBKD6LqX95/Z9tzyX+GZx6LfwzS7+4dzIkvKJ9Ma9iJH9+kiNvl5zd8APo
dDxe0wUARkuTRm/48C8uKlKQrW2r492HsACjuoUXbErZatuN8caQTsiCaDnT7CZ613Uyg2XKpZM1
DQy7OfMZNS0bMPkcySi/z2xIP7K4Z2jVXIhBe4dkRoJRUZKFZamhTu1yXPbkyeOABwIrjkCxcIg2
8hgoTIsF5Ez8byKIKm/6AkSiEA2PtbCeLDjihOyZd3TrnkgoJ9IPa5fv1pgpwi/S5TcfL5AlRXvB
GG+l51RrLPLkw2mT8y2GyiF6wmKUchtfi/GlVVYF04bUQT/TFCzPmZWSsZ2zcPdBC5D3uLXe2ZZg
Lg9LBxuPB6bicubUYaLNpRIqL/L4tVoBaMXnmvGg2LqEhBiQI8+0d+HE8oh75cg58EOYi+ga1pXZ
+PXhxidwMU9dYMmdVzqabKjbEw5albrzD2FA+dWBldS+1PwnP+UoicC31zd7VxajlaUk5R6wyPJs
Oq8ZbzpczsTAux9+hg6XQ8+1WNOkrBKA55d7Zo/DN9xWZoXGzmm6MYt5HdeT8GIfxle15YaE9zOO
1D+IYsa+VDeJiCJXTiGtu9BNOG4kTpdE8bP0JeoETQBESs+3MHM7rxWUiyLR7344O/JsOlKjPrWS
SXeZKuZTCSGRIxPgYC0DH0SqZTSc8R1YckG6mlOvVGZia71Itpty20mhWvDU/vOvRA5Yfm3DWcVH
/xFSmnEa5J72w1yHy92BkD5Ni+D4Y2SYtmUtCVK2pOOTebw79ODYVnloD2bmNLqxJ0xCf2uZTiXj
bgW2Uhdlv+z4SBs3saQigPNsrPXciVstYH0oukAvDZT6gakdojtkuJs3O5o7pcAFwyWlVjrsZXnH
TGGCAL+Nu9qcHu0HbJXKeVQzWzJw0jKfMYBOLNp/kc9c2EdwKKx0VttuVV5+eP9g30EVls9chNEf
hh0R7G7V7mXxP/EF7z3JatGvJcS3qDepNcpc1fUI8hdpYqAaboR/PAdz98IlF5XW2gUlSYfIH8JF
70fXoCjRGJpzZYgeoEFs120iQwy1AtbXPubJJSG3NRvuMyQXKsIQRylyQPxrGa4t5elQsuaZXlWW
C712NYNjGZpTc3+ZYGrHFTAeqlrI1dz6JD7vK25Nc7b4av7al0rwYrh1cndP72cSPeDnVfotTpMi
QSAap9p71qTR/X+T6LJjaRzO0ivM/L/8XyYBQ5pQ0YLNSgNvXOfW0BUByhzzgbZjXgU3kq+mEpTf
LsAmY4yOfANbXCZeDng2/Gcv0ctOaeGDC16BLdgmkZtbMwjLbFh/MGdzQ5Y0HXezR5+5Vz163D/f
mHrqLqzYC0WJVXS/+ALgBFdV3rcM4w526HglOGUkYtTniBJJaaS7phhAiv6NnupR4w9eSdU6tcEC
8++FLBhEMPfvN0W4ApC513JpAUX4l8ROsfVwtzzuPLPZdcXpvECfyOj4oEsTEzTHMeRcHyqfWiV5
fx/WxrIJU92p7Deji301IK7a8auAHcaOshK4FDST+3mUN5R2gquGoe/FfbTFX3ttziKvhJiXoUEA
P8jmgx0/+9QWwEauPCyvcPqa0i4q8g4CPKZgj9QMJ84mTk/zJRvbpJ/4/KjUjP/MwlEV1RaVRf9S
xgPVAWq4Ls4AhRRXpilB8pYni0vPXS4vuAC1nyGE/sc9vXgqYCbsknFyR8TbE4kNNasZaL6k4hd+
IhNAzM+OxhrdGQTZMagqaTBT28wOFfSYJC34UNT7BvAUD2iw0QFYAlY3mMyMndLtiet9JGpx+Cou
sRGLC+D1hR5OdAszOxRlJfEnxXFYoFX6LnFYP1iOgLIHooh6XZzMa+UHcfQWnBPKHFgpgT5IMmmY
k5PDUnDTDG2bX/ozcdiTjfKGRFWVZU+s6877gNzttRF00VOSVfFONl7atRWcdHpqmyQxJ3wtnHmj
80VnjZF9i3XTMNxmCTXi/uJ95KiO+gAU0Ye4gZ9B5t/lOZWD0nAs2kbrbkLCLbfbBIKim1Kv9ktm
91xGNOxKkpKnvsF3FCWQ7DyYijUeW1dVejJ/eC7p0D/GS5rvUzLsMMpmrk8c1K/oCfJNQ7oAOxvg
8P31tKtK3p8Hd4iKLcLoW5laAm+T426I61rYLu4lcsnkFk0gLsdXs9e0ff/ZjzOCIG8MijBQKcF+
cYmpDuZdxbf5YNUnWH/3ahkJAPi17KcP2B1XEnwxlBmr04ZinrT/e6Z0ZjmQ7d73PopLV6CiwBXR
5VTgbNlN6fidLlZWbhzsUiakJ0pMXmLfBIj0og0y+uSMNh4bmD3l4kAM6UhLtn9mVR8p88kc4Q9k
Uc5uFM4aNRwF+sSXKjwxMmtO/qWsAPTAlZtFK0wG2+yfD7OardqsXTTQlDG8zDra+UCuWrW2UWOG
zxDxpefh8AoKDMg+of1G+VOtOGIO3Fe2Ps2z1GMg5iO596YFIx6RLF5It5Po9Crvx6XSe3XKMJx9
SaYPUIfYOZyL4Evp2OY7JkAmp0d4pSdWtYHDiCe+7STtmKmJeyxaxWe+hITvsI0uBJPkr/IC5qXQ
aq2q1ksNJe57PXOL7FLW2wtFTbV+OGwoRbeIzHulGxvk/cL4/+qUYpIF+xAP2mwNK8tmKGHqztxq
Xu6PuUgct3qOF2FlULYnVynZt+oK07g1BwKnYC5Elbfp3WogBIelIvLlkzoKYv7mazvHDVfotw1t
FZqHDK7JwJ5xpWfkk+ZrU2c8/NGeHPTDSs4M6nNFRDZl2xMChXGy3+JuF1EgMrLZYDqYM9WGwnMH
Errdd7KcIg8zuWlH9K+tu6LmE8uEXLPJw9SKohxuspNghgLcuXxriKnlwjx+zlT1wtY2jJqxXT6i
+bbPyPF4z4FoTgltKRZ/8HellqiHnB24fxFDyDfx0Mk4x8HWDyhxpjsbl/d4mZHZVbotovhBEaGS
9VyIsHyHfyqEZnnCy1s+WRof5LOeUdkUMo/0TmFZ08/WKolVLU+Kzh2nwLH2liEcZcYACS5Wa/qw
lLYqhobptyPeXDPyG0oBefDtBD5dZW4+QA9vHHsn2yk1ZGCNhDeFDtWK1toyKXwNNi2H8lkVBFBO
N4rOv+F/Ta31WoGUpLDyJxnlX2ZaXBK0FrRo1b077UeAX7ozHwXKeZ93D1HdDs8GYFShSvKdb9B7
SeKTCqX6aebqes5B1A/RAfemzPOzew+c2XWcF36brqyTIU1SNEOL0WLh+1EYK/dvusU7EdqJuZfo
jdMLsdr8IIXNAFLAxzkt4618ruaK+rWwNWQ2+ryTuXGQe2bReF/4gf72VjsOk2XIO8Yvfi961S6x
y3Eqtbj9gIL2YmRguqtJpiA9RSJOfAh9ASNBzf1YABKnzEiLQe44rSGr3u9O2B5qxrtR+jV5eagt
2SIoL6E4xQHWtlhAd1eJ8zJXDm7lZ2TEs2CIxO93dRN6rILL7GlaII/VsHE4xL7gJLbxtKMsCXyv
tCNmvWrxQALvajFdO0PVzz0TBP5TnT491lqJBMXjusgKLJCBTCkMfY8tDPZ/UYNME0Qb5w7u9Jik
fUmr3PjYo9oPpfC4ho9Lw3Go8wkauUiw+NGPS1Y8ziQm4GeRoCcCEfwzb03FPDdre7Dixy09nGTe
BwjoLzhzhie0R64rymSqGBKZogipja5eGR4v8KeOgG4LX8OiCeT7AXTQfRu5qC1cWyxvjdzn5dVQ
BbCUKWCptIiujExmhByolHsBzIuhGt5zx9+LghOv00JP7jlH8vHP4fNCSbgwDARUwjkXO8ctwtAp
iAq5aPu84FPwwAkud1qd3vZE/vFrYJFMRgvD4+7GL2JTy+uTixEQJciqdlMn7BtmWlKiSg54zfbQ
FInv9e7z1K/DqTPePBAhlrA0ESCDa5gpCpmVluId44oMvnHppIhmA2XQ3hmhuz2JdljBZcMseD7x
U5coJgeK0yWpSAaRL4P46SNXCEbK3sa+xNlN7riV01snUOLgfIIo3F0fl7BOp6LRgqM7xQchqopi
uKIas5WGPqWVDvz7x7LUlTvk5WUDsE+J3QfnBaNX5ZhxGA+C8dl4bLbPnGvadGrhqH12GfVp+MMx
69CCWMG/Nbq569PxgmQpScO/z7zibZGEsylPAZuZFfQOFzqfG41QUAPlxMli8VgMpDMELNtJwHSa
WW++FC1HgMw8+GSQVZKR9SjLFixAdeozEXkC4uHGvREqWSBYzHEOoogOBAcryCODLNU7m+QAmExs
D/6CrZqFDsuugXK/6cAMJoCsoYvzWwJmtAl75GDohCvPL/vDW81EqTi/TqoW9FN2whaRlm3PqTHL
2BGSPNKTNo8vtFZWsefCc2ypsFekksEHc9ibDfczMH1Jc1egx25Bj9fWn/qyhjRGzYScFucU2K9b
/vdMA9d3PrheJXnzbUs/xiCEVx+W+Toswj0wrBDmzU74OBgvT0MJJbU0+1xjgsO4jE8Ql/6W+1+K
Y2UK4b726/J1JgGFJefGMrsN7xDidtdXo7nwE+e5HugUfQ+PagO6oTZTprpkXri2fInPYuQUaXh3
Zyvt+BjBZzYad4oHSMvZHOtQKyEEicXbswX35OQJrLFDSeHfoy4Uf5lJygRbiz6lgQoyv8jceSf4
Hd6cIP+0wyvfBvGlD9KGX0fbX5umChHjlv6CoQ+bSD4A3zBoufCHd9fLUFC9JI687vgBBZ0obthR
DR42YOAYXUm0GylBXaNRk+UQe+bAktvSXV0wahRbLPnPxGronAZFJuJ/WEZGaRAM3yFuiKXFnFi+
ci2xmov72WA0/wgok6OXS0GuWyhPFl0cD+pjH458YsYFu4e6PvRwELgbf7dPVm70ASxQUI9OKpZ8
Iyt+qpgWa6yUyjy7V7Ql/7+qqW41I9JjWRVae0YlYn39RMPjf+QhbKVmicGvhI3HxmhzrJwNxOQV
cs3mYK7W+HluM0HnjtZb1yMqzHRqDOfasE9U9+LfY+yAfcSKd2pL+IboxuLxqe6CiMaYaSJ5eXIS
UKNvbBvjoWYFmfHCCkG/jQlwftpXDz92ye6nF5kSLP4/hSbLEqDAVDwu0H1i8xavJhHKLFy+UeFa
CXGPPlYkFaa8iRt9rry2Rsdw4ZkayN+dEysYGOOR4URTG8d9xa4Q3FWRKhOgD5eGOGcEb082g4p7
/Ct4bWnlFmkjp0fhq+BTHzWS50+QhSK6BP3WxpmkA+MX3zIfA30EiLgs8yrmoZdgFbAhAZdteAWM
IPuvqAlMcgAKJdJmQx26ExGG5F35l0Net+qWZXu4zwuEWuYhKrnteIQO2a8GmgzWE/Mw+xpdDz43
FHvn63ycTnrCSUaMy6pEyxksx86RXERn8lPUUYTkcU7a3Zc1jRHD5R3Nl/zyXT1ZN0Y76hpTIZWq
I315DzXddYAgHmF6spVfxPUpopcjKQiMLBLm5xzUP0qSVp5HAA+tbBqnd2v4uA51IKrWiDNGnc2H
VpAFhgQVtiCQUonSUwARbO959anhBV4WZpJ1kncDzpbKCQNAABzsTyrmNBYfdoUgIPEjHWpl7/5a
rvmqdjTN9NY/bZS5yF0JhTYmSdoHeRo/xQIjMHgzjE2CdVXpon8csys6afyJZ9yhwc6C6vmfSe8H
wmj/fow9wjiy55eiYLzvz2D0DWt4qeNG85wnSsBIciQ9peTfwL1lhdeIdhmNX409WB2aJ3BkNyEc
KYT6+LyGkoq66rc71lrjej0MQkrEFJ8HJQG+r1nINeERzzigoXEvkj6ShrA7NN3h+zeHGp0mASZm
VHPi27lI6NKsgclwavn4OEgj0qPvN51lEdm/dAscnR0a5P9SmNLKfWY9FoniZQi0i3WVc3PQ5/it
5cPfWTETp3QhuutuKdlfnAGqb71DD2uhSonUgjT823K2h9hFayqFjG8hQZt1r1sS2ZtKeSg7QJ8Y
MRVpL+5qG3jbnppy+JkSLQIabDwIWEDX/quSFq+AG0Z2cNkzk4C8ua95kmAS1AMly783pTxZXDTY
HFpb3IovwSxb/+nHw5+rus70HQpgZY8u24sWUvUctw1Z/pSYOGXMw7ZLKfPSe219j5L/vpGjkEtM
6nDL80vfPernk3A47L97aW2y8lxpdj101C7ihF8F5y8YUO56qdMqMoaFMjkWcQzAqzs7FtzQIcqU
xoiVUESPM34TO6Hot7MCHE4BIa96P8CgA4Gi24o70i+JwIFJ5alnOWzx51m8ZpRhqTnHNCaRavNv
DuyEWhw9VXvk19IJcjJOdIveajyKlB1iiYDUDj16ylK9ZUiTaL9W1OWxs92MveaPQLBZ/ETC8d38
tpxCa07mSSfzFK66tEwVJjSirR8LRK6RJsBhqq6uoDDvhbDihTlQtPulPp/lHMDghLE3ZO0sa8s5
dbTVrvngMqxO2In1xfQOjxkOXT6wLHtT3M/IIGEMjWcGqvdR7y+vqGtCnVE9w2zmsBpLQ2hpBduN
YTEOZ2obSXz69u2p7OMefQmD8+4q0aj5W/QPT7T47saD8j1XvOd8K8oFvBOFa/W/qUZnSwxV3MY9
iRAoKCUd28A/xQEf80zffbGfRJP4Jh8km7/1RKePwYoDGNKYiJrD7PGuB5xJLSO3TS/EtELatUSq
lsSFYqIrpjxx2YViZQ+xJojOxR0q08rhrAQTV0sV2gzfLotO9TMbz5s1wQIPSlIx7z0/E967ojll
AN1sA2CQOB7gNKqZLeK6S9VE6Fdu/C0VnJsMFVxzp9cDSgCce1S0EgLf0RAzUXEDCuHDX3lZa3Pu
jOHET4+Bdse7dD3iAuX7C3O+3IRlOVVzsJopf292fiF99L/irugGiQy6FYMB1w1KLRrRfltUcWrP
kYWJhQpB5t8N9KpbN83H42Ipb67uXgvIL8D8eS40A6M7uRC9RF+BmrX7WPeSe/BCOT8Vyyqpz+JQ
VYJEKkBFNw2IoxKGXWR5xdyKZ5UV+zcQQpcFMJFwbphWRbOjFSVAcjs5wQiQTESlEN//PGAeYg29
SmtjOXEjjeDerAARsYcOm9QfbuzQr0J/XtqJXPbR7+2NNxChmc+NEl8ZG1gV+dAoGubZ+MjcE7Wm
V6mvZxIfF8PP/nFSZJnDutc02gJCQd9KSLFVYhHc3n6V9fDg30OKrJW6+q1p0ZPJ01rcC/K0gPol
8DgabXmC1yQY/6s6Dc/3+dka8oIQubLh/OTJEiRTjRqiDIXXrgcja3PtzBvs7isEXSdSs3aKiFpj
8jNvQcgVByu9skDXnLqe5vv+r/HQ+0AfbRaZO0AZUT/w9uS7JQB58jNmAGKtXzLP0uriwqmK+gsK
i3T7zEfsyYr2OFPwOcmJvKodkCCpxttnHqhM1bLAbmkqB/28fQ/UkCdX1FhQZHkD3S3/LXRLrWis
+eBEj5bFGs1algr1gSMsn3i0T4WD7PtD528gNgtcfp7WpDkcMQFKnyqQdDWKJMRRotI0KYPZpx/m
NzF9ckoZxiWZRWd+CIFz/FTg+urvFQI/cE7EQcw9VnrbNA8FrPTktfsZuek+DKO30GKl69gFsFKH
tLZi53eSu0Unva12vkauPhz1dws7yMhycvOmFhcECCS560Ntml+dv6hXN39A3HYMRj4smf43yqWJ
T+Hvmee0v8GcC957hc3VrfkJkQXWtnG4QoUWqrfItw1c6rUikMhm1bh44fUjX54l7pwa4l94jjMn
iXSLjR/4zVi2OEDu558kjINqL3ywHWQVXBUY9uE+FtRPLYkpxm5DOgFJIvitiQ4RZHGHZ3iOtO8V
kUK4k5D68uceCQY/q9RdBJXqhR4vo8ps+VLPY1iioLqFpMvgAym97e7FAWdq+tiFiZ1Gcp69sorl
AnEX/nsX1dzWLHVXJ3qaBY2uJgl4RmMQNbdkAJm89XihYGx30wt7ZdnFwOXkNeWHwypVZgFVSWkA
1w2wANxe7z+WaVRkrQ6+SMfwuVI095bf2LRo+jiHg/PB5b3gfuTu65Lsgu8H8/tKJMDl6uJr1ZJb
U/ZkGfXTw7yHKWMph8tO4dOoPKBLh9wFR6E0T5SpFifNyWLIDCgTS0RPo83tGcxa0cIk4zUUSgyO
b6G5RyxzEBf9/8tNVA3ru+wGB0liWehPRuE6siLMtfCKPp9mEmEXsnORl9TBQuHLq/akSBuuapb7
j8WL4IwMpU818B3/uZSGjEmrLhf2qUHMowXfTmzfzGuoMdmXW0VekDbNpkoPZZB4diXU/5OlixaH
z95sqrPT0EyJUuv0gOlpS2+2HKtXO6+RmNjZN/qQa/pI4lEfg+a6nbvaKoaWRQWCdCaoz9bL14oN
fNU6H/S1r25L3BPT0xKsxYKw6MeNHeAObH55Rp/wx8ExCRGqZWfeKUrapt7KFeFZv2NnK4fxETCF
J3lg8fZ8gd+1/xUAj/+oOmRiYKlPQbCi9WmErgdGfmxG9XnUlISpgOErVeIakf3hhy4uOZNpSi74
I8JgYDwnZj5WITYxHEv5vafiHxqU5DmMSxx1eC9p4YiNT4XdYtSAIm8lzuGsNRw5UMkd/gPbVIKF
KjrV2tFFxPrnTsHjdynDERJj+opcBCSK1mwCtg3HSk5IN+MReVRkm4VNmvs8oKStzo7MpgKNJMpM
sfTkdZVLew8PaS0que2SdBhfABy0vE31DqZu3oMlrqG8J+kugGml9WynxWFsa0D8pDDM0y6HyhnY
jjXFMIZnuF7uuUGY5aDxrszd1PNJY0S6Cj7chCY/xOiV9waSRLRG9OuCs7HcLjy22AI4adzehkzh
BI5du5FcaGg6BVKm4kUuJ9jbpnKpyeIAd5P7rOOLAfd9TsY10dVp45zfTCaMe3TmAcE35MsG0X1V
pNfhmAB6HdiolBaBY7xBzWOapDJ/ga8z/LLwsqya0pZ6Suyjy0UG/Xnu1yEPVBOW8EW+eykVMeO5
2n1EmJxqoBUqU0rL9D5tw8rPuDCNxGksogtoZYlWYKYghwZj31C3w5fWKJTQqm2md4i+ag9XYO90
sL9Grba4ivgy/9ypfWjDPYrEWUOdfxCjTSingBFdKlBsdTa4XNtqq6gEGlHIqudsGFzwSJi9CYak
XCMmjfkq6fHJ2S7k5G1Z64rGpZEc4B3NNWQKya7sttZ67APtFxN/u9riKODVVSsPnzNZYcxmiY8/
CoElFvyWvwdJGoFvOghLEYXJXOonzbJYd0HIYCDgDfNuch111lhEYgY+SALsJspTh+7sg50Z6Hl6
aOencmefGXm+t9KN4Qp7DyF2+A9eUYjbL3GPbfzSgUV5aF7JDM7ZC8YP26Q8Jxf4fP+wRsMkzLAo
7mR+VAn6xmI5aYY3NtNE/5svJ0Mc9jDHS8owGWArIB7KgpUPLcO92jkI2xRn2HReUHU8IxVEwwuF
DelRZWZQz6XQZzRGRfM2dznp9N15KtC5aXgml6e7I0IiAznRahuOQokmx+UMtRMzm9XbrrxyMhOm
OYnhEJXwWLp+KYAgUTkLCMgpsShlud5UKKTH9fi+HgQFPpvbbEQkCllxgrTBEaL4juDtt3F/zBTe
j5JPTeqOl1HFmMxgtx37nVErOQIHIR1ONP0uVbG4IsFmG+sEJron8ZNrPwVFnn5wadmch9tJ5Yju
A+CnrG7P1vnOGDHr381+OGOZuU+f775l8nvHQhDxkZopgox+u4hY6Bz+GtRHE6iekdyk9+wiZ/CZ
hxELAoJF8FmvgQ5gGkezkqzEQkv9SuhrNUigEtdTKLIMNDb+YqhrZ9IPYxcX+++2tsmbzjk2xiIr
8LnrjDzV6HhfBYG6wlI9+xarStkdrUo12jNyNwfeqjHX152s432CSAigehV+0B94mNQLgJUKu+oL
r1KxyG6+rD1sCi/XFELVdjul0NiocbxdMKZk07n7ppRojt/kwel3DKyzjAJGO/f7m8AhL1uUQU7f
Gm20QPm+7Y7jQndbuPbUq8QDk4+rfhyPZN5+49o8z5u6us9IlvMb2lz6zlQZ1VcdvmQILD0UtWv4
Jw1bdxYV5gExz/f2aWAQb/dsyHJexm76khxNCJvM5FvihcucOBJq3MkBv1GKZlty1TL6jpEBEEJA
ShCr0iRJ+uy0A2DjqwYb5LJjDuUX+GaS2xu2S9yrax7FCEnOzV+zbB3WRoSQSCUO8WpafRH4uCH7
dw2iBUw9Sabxwas4eCfvcmYObfypWFBOysncQFoSXrz6sROVpPSBg1qn9HrPt/ZxAT4f790GQOv+
iiYwW461wmGvi09DwOzv3AGDRathU1QLI0xx+GG89frWeb0mrzZs02j0zWCOyHZdVHYnqKZhbe21
yUFmQE/FvYYmNuiua8aECT637jN9pg2eqp8UyqdyqMAShj3NBrhUJdYvXFOcIj73QYZp6RTDaQe6
K0IvZQWT3hD7y/8Jt6JX4zaRph0sJOtxMqZIfuNzojyzvZ+ttkUhP13+PpALKKtFWJKLQls0CgQ9
//zhN3wIdevHqhBTu9k9m8eTvo3pRVXqnNx355XlS+m44U4FSjPNfo7amGbhx6Q3N6RTuXb0nyDP
kiHFKfZpw0usPqlEchMzD5Qm7SGGQOU5KbG0T1iMcJt1RrdoZtMRIOwWYSqvJQ2w4Cof8IOhIrNR
3+EM02ynr2CX41EVZgaYmb5tj4b5ngjjFbQEqtJIRHPM+1Ff4R/9z2GcYmijHdfSugvW+3/0Fn6e
yX46Xf2XSsKsGYdPDYK97cDkGFFVVZEor7G6JymTX4SchI1te3Oz+dvZ6yDwrU0ruqs7V9VVaSWn
27Lq+9Sd+/zJ+7Q7noGiMTHbqGaHpYReP2QY30MZGrnwztHCSg0nLeOXLowxrkKVl/ZaxDft64Ua
DhNRd/wtRXkzwWcGYGKiXbMjrw43fFImCK6XyF93ypw4OGn8fFAivgX4l5RJ083XHT51mX4DzXOk
RCnFPF7zvXArPTPf/7l03VRQ5KX5/Fia5b89aKc2sR5Afh8rAkIlD61jISdFAI2mH0Ru7Y25t9UA
Tkd4zde7zLfqDOWJOr6Hf0fxxVkiFVNzudkv5JMxPe2GXBgLAMazFPCTwX+0q4NlEa0TNrea5y0Z
tnwbe4T8HaaNxB5GzDgNbt9O87dmr4PsjWiiaojVMfvlb71ZNfa4OQ/qUng/rZ9b0NjHidNbyWvZ
LIanDQgfA/KMDIOg0M6RBb8aGaQLLOxkOWHX8eJeW/xWb36rSQ4TYXJMD4i3HseLY97tGtMDTQzK
V/jOxxOMoKN1t3YEcYjwvcOXxoDrfnmAdjFfNfR8jAI7ivbuUAQakNrvbe13mbw6fC8O05wMzD+e
/eQLH8p4eOpY+bIfdKikgepKhokzsdjsSwiimeT7+YMhQoyEe4zxHitzyMjG0S5JttbQtMmr/nng
zyA4Bu7FI02IvTeUxsrDu5nwSorOWAyaZcCMvBt85PYJGwPeXX47Q5Jz6/69JKbjcaHm45uFrXgS
2AUhOA0AZA9H0WWis6JmeIJBSH4J7zIzO4KDsjzoQOW8gOnXjGxU7xLIpavygc2yUd900KnInElX
wiQyAjyQHRCqmGJDoC9NHOfrAkzpt5sL8O1YIDhGZcUXi//HysjX7rGvJUcGMd2Mdlkl1tYYQ5a+
j2WCu5jmbUYjnQyI3vTv+l3fFcxNM8+RLCSWkxwzw4ST1hzpsRa9DK+TgtCYd9bbIs3bcza4KQZH
eOnurlCodfsC4MqEUDQi7eJclpBxjokL/NXhY6LoNLEObQJ01ScsLmaQ0NfH8AYNIcD1oVaWmc9p
PWVoWWp2jfDPu8Uq+bR4pPsvk94a8W0JZQkxOAvywa2IYIPrFtxTlVhS+2+sDFx07McRJ3g10N9j
2dIXjxGnP2GLYlWnjwqNJkbEImb3rafy9QJZFi/URrLxjYF+QAMtYRDrnTEvUaL5OF2uYg+TTf5y
Jb0GaPYYGB5bdYgoP2vmCO346rvpMUb7QgsjSbDqvR0PdTpe9n4E7h41evLtl1MKfQMU2BH8HGWK
KdcSnOstLITVd9OITLH8seZDASdGA61hQFpQzvvXamZTCA1/n1HpBxT4WtO1W3PvRaLwR/FqJ/JF
dhrSl3D6GbIEa/3FDEV/L74MD56/VYjWJsJrrnIdrDNJBR0LEl2n/e7w/2GxDfemzi78shwqFfNa
AsAWqnR+QWe3gEoW5AnkEve76st892ZTOpuyc0CpMJFis318lEoCAsr1rp1Zm47WdEbVF73RER13
9rJQO7n9Ahq6quxgeUAFpOkUDw1+uI4xzskf6ByVIC7vUvqR1twNksWuAjx1xeQFVUfjOr3GuBh+
DPJG3Ekb2SQ2X5ldgoXdv11f0nPQwEBEJ8WwTJBy0TRZKdDBjOar3IGXbKEdcp0Do/d5MSuLbPPf
ggOI6ymydb760xcpeRdERf2ttBu01M9A/gfgs/X1GDF/5Yq3g/fJRlvsHNq6P/pfeczfPgY3zNKR
ufRwcvR0Y/iu/TAC3s1nt0XR4HMI1gWHbNOMbRTcTgyATV9u6zrKj+fb01YntjpDQEC58FSJ7CmN
iPrSYmTs6MwUwT9lIEGe8TOLdjerbGo3gVNXuKFj0qkOZKo7S4QC8jf4sfs29ItnySrhyJp+uRRd
I7Ah7iapt1cD+n6SfvR310u3dQHF5mZxqNhYhNEnRsqPoy75thvFqvgS7Zi7sr+yj35ThLimxM37
zKmNIVUB6uSEZEFwfsA5k90EVG3WWbdwtzBebBxGmivGVlonpFfGWxYWuFunszplKrJfv72tTWLQ
ayq6/gwUAxbHxufXJD/5FqV4lBVxa/JuKNPJ73iR28YD1xNLXPc5N+1jLMNDhQ6GhMCk3D7RlEo1
KPnZ7i88gbWWQClQyvt3mY4dOfO/SURjJ4m9jE+B1bcQPrssFoTxdUiCja5rGnWq0D7hLRS31LAG
ug/Giy3CcpvQfRfagYiPSMQgLtV1abLl3uIr0nrAZmBqZd2l1VJX+BUeS+qHNBu5PkOSE5eLDgi+
T2FrSr/RhVAbkfgIHAvHUCjsugWRvIE8KWGELQ13RO0s4foFXnZZTVETr/yDhAXCgG0TJQQyk510
tutpgesA737AwoeBaNw60KxWPD6GVe3XsJmerv0fOSAaaziytd6WofF4MljYe9GhMnpLt7BStIjM
T3Jd8+1En6Qd3IqOU+qF9XE1f2XHqCOVYsJxBvHMT+4OdR88iCvvaWGvresWu7kUf3GjIswU6y7t
ZFKmOj276Ar5PthIyt5/IKqOIZKGlTl3dDFVO9Ni4uR+mMmWVGZfZYZoBLSohUTtS+E4p4H5LfVo
sbnuNz1qx9gkM67R/mQ793a31tUECy6KLMiZ0f2x9Um3NizBvNO3TFMyCSx/ugMoUxWTovmssiGS
xj80pqmxQ4ba2iVFNgnmO96fJ5Pfsd+Q2scZWAobipGWyLqf/zvjdPwDi9NHjavaKkwuyEPoBVTe
Ek9PmxTKGpRDurtBnmG0qRqdIPZ1MxaGNW2BiGEl5HJCM7w7arRveqLWNU2R/e6Js7H80HECLGVV
dfKKVP/NOQhEZdOz4MElgL2VRuUdxnVZ9GDrVDw9z0q85ufYds0HF2lj5C7E4d/gi/MVuG++ZnKs
DG1+5UtR07vq60aO2+ItTmuDXVY9PmM91Eg1xFLatEPy3VPUcMrRZd+uGbeoY+unTTduxNB1IaYJ
0Tj4rupDOdLIineg5yREacVeQvnrTbxepXP+iIT0/fqdu90CQm0KUVIGGJLRS2UkH7b7SO9CUTIa
zyNeCSo4pv4ovwHQmaI0+neDt9SyjvR8NNf65xqSlmtXnRTx2q6WINO5cUUiVpBIR17aoc6DleW8
AeX0f9oWEgObdLVhuXfb1hwonKck1NSWxdpPKY/m5EAIUDhCfKxSIz6O54GdU21lS4mJq1vf86f9
g87Kqte2Ic08/Z3znw44csGGDwqg7elsIuR91ja2Kb9+CwYsOjVaH54ao7QXJZKp0SBcFg3Lp0B/
aBN+Xitu1dosRvgLW6xjntnNDJFScijZYI7rXuET7EBFhVDl3pr+Bcvo+5Pm4klbpEFkVGkctBoR
rM5opcvy1g1TKLwik2Hka1BMR9mriwnMXAsdfmofxoFa7zXgiyL3ZF8/Nfbx2fJ04rDE4EY0JNrO
8MFy9POG0bvbPcA5oGNQQTELfmV5RvTH6A50kouCIZLJa1XuBIgsUacFwyrAlFRqSHtTAYK/1pUa
K7GtwDaqMq7A0TZBv+PBvsNbrfLXSIEneaLIT05VWr4WDdgYdp0EfSvVEC2fU1mw2TbYjpCIEn5o
1HSQ5U6OqRXre/8ISLskjVSA5UW7gmSuF8KJGtZm+l4qVzIyrfN5WwmjLxiaUikL24iI628aHpvh
PLuQGRO39WLusslKBAzsq3s1sENhEsSZ/7qiKEnSQALfytxENG4KXfiUAui/oOLjjfbv0YsH53z+
dVYsxyesribJHYRcus1vn4QGc5rzYDa1xsIKYxsxcv+XT3f9vo8lNtqie415nabI+qxv2YasvdIZ
72fqE+jThz1/WPlf3SKeEuSsHZjxH4v+IJkdIe6QJZBGyaeW1xo/q8G9vnXV9O9v1tWLywzf6AfY
6WRowkvs+HxNajF2O6zlKj3dahXXWvUWedHvOfXofOSoKtXgkJZBkXffX/Uuj09kRb9sPetEpdS6
cjEDOc8+4vFQx+Bt6ijR2p193k3zqMlrUAAvhR900mmvcTbfXLgxGdJEyvEvIl02KvMfG3DXvOKJ
FWHDkiIhEGNJoZ3bp1BSw5AnN8ePzoLCzIvNBfv64Z3shOwM7NVvRoWV6tyxeXDtVmFMvAGvkyDw
Bk9jKmBVycrZ7XVYUMxXih45h11E2rvNuBuYKLkncRWYKm3AwWsBygcpWqeQgV7DIOH8EWxmS471
X3N1PVJsTVX2dqNxhvhYsv1xfx4jQbHGLPjGlboFuN/hUz6P+1w4C4JMq5XJdSiHRKYnQdmg7MVL
I0cIOCiLQcAXT9nM0dWLdCt4sXuUdlZmQpe2rLedxd23GITkIL0qTVeziO0ndcQ0DqdKiyetyZHE
sJPQLC+rW83dqnLZTZwVFciaX6TfCQPD8DyKy9nPOScvcFAHPAxjc6Nrto2Dhhf7Rnv6rIwrhw9B
HOFNI7vXAdcsfFu2G4zEIRBwtkGOYD2k8sTNooWP1YzZ+snekfgAQpZPAeTGrdrQMd2nywOVUxXy
8YD6teNE+SkT987q+dbT0YGM89eb91/Dpu29uluH0NOUdq6BfARt8HX0MAzCgVyjzrMEF0ybWwMg
/fYs9zoxJxpz+wGvZEvmyXYRHiUvG/++65Uv6yPOuTezl2EyDGnVGnKu7SRrUqvoibDSbp3rZz7U
EhB0doWCNdFn2SGNdwjWXBRXAJUuNpN0XegxYE+iVfmKhh69XgiLb4M4ETNNUK8fScZdGXPDT6HQ
9OrCGQ0ZnycNlIUXZ1umwpFLd6j7nNui2JEbS3YvqVXj4+zo8nthBINpvL6agiRP+6P7S679/HMM
kZ/GVryTdP3F/sUWQx1mwYoGhhK6KX6NqqSN6vemWD4DhANx6X1ww/hTjTC3W2i5L2V2TtIg0Z/2
+biv7ONFknoJNiBkmBmDkoJQT5MXOh+B/3x8jMJbQP+vVjwOOGTQ1H6gSDlniP9v/7vnV9pNJJzu
jc/ngD3q1tvu1cQ6yRrEftautvHSosAewYoLepbqWDzR3V/1c5c4Nw/+Zwso9nsFqO/+vd6BC+9G
V5o5SOMZwQgAvYcUNkZeLWLBqYy2ZgZMWRkuoLRxTWnRvnbIuoHieZv1h/oAKD9qLciwoRgkDuxT
g7jgv2kGsJlI/OS7rmCl4zqrojHpOK13DRE8w9tcpALoMSXerB2KFz4gPzKeSz71qaeXooW20V3n
148H+fq3MT41YsTeQDZ1PUI+PQEvEMCDImpd+C5REFMX6IiwbkFvNEV9GfWqh4oF2QhmXwzOAbP9
fb+bLCN50OF0MXpC/lo28dtttaoKZwaVTZ5UDRlRpuYEB8/tHr7P8ZBHmKS/J3CN5H0ZgEsvo89F
0AvIGlPX11JaY8LLtTJQ4y1eKDfRjf7JnzgxIjXeoNyf59/UUe/mmXf5ng0ZX7x8d4BvryLb4px6
/5xyhErWS0mgqpBFeyWq2w6OOXfHYg1zCGKrFyg36zYI5k+MNxfF3+4UAlZqxo1FxYdVhtrd6Dii
G2V9u8qdcrlgA6hT6ToiXEpW58oM08zBZ8aiARMXEirjZst3ZgTqHdwdzlLwI76MjVYH2WBE84zp
KqxAoxBUt7mjHgHUVL6sNGVNoCBdwdIQLU5VxQzWLpytl6gbbwtp0nfbKMADM9VA5FmStX7OUzoS
FxgWztNS04GtDkdue2bD1OiYfkMB2/m4gx7uWIgBGDmxEmqrWLmvxfbLrlMNKcWhCXFNAvFPBgF7
Bv0V8h0v0inUeSYs/rMbgbmekXVgTFISvVLhv0fvQzwJrfKw3BjpAmTfwNdH5s0ENV/J6DnAaFYD
WCYRazIEvkGsyP2BbR+8nROK9jj+qhrR9xMr1KqlSIwzeRtG/QeSmBsE3uBIjz6cIkRN6uCw2kO/
VsNNwsQjmMgK8NFqbnzohtoHyjYt0ugLzVDnBm/j7+PlX0kXwcqA2pUF4NKtYKd4Io9IHgTKOFEE
FiJyc/ZMUfJ+z13MikJFN74dl11HTAXNXdHKLA1aEmTM9cxJQ8Fj+aGD0h0ARjQJ+j570mBt+eiI
x+fOHBPTALUA3Y2vHr6tEPRTsT4t4jYphE9TbvT+FLCUHTJFKhzp3gN1E/O6OG1Qp1xFdQ+2Yr94
F1CmLLkCHUDx24mGJovHzaOioF9OzvVVtxEtd3rqBUK22+OzNuhT4SiUNc1PYOAlCxtBzk2AwGc0
/6MuC3qd7O7UiYOtGSI4Jf+vnrFfWHZn9b5NNG6hUiW1JMUIp0vRhgDHEe0ljTg7WUFI3b7TxDGP
fmKRtjQUCoaNEmkI/aGdyhPIJxyGoA1FRnZMydiQxwnNvtchIAOCBdOYeoGXtMnDJGC2gmiv61bv
p7/6uhBefa0/e+ERVlWXU9MecXZcUj6TNQ2pn24CShEawg2fV5R5GTfBFimCzmr8R/CMnSAhdOuL
8wbvOp7gLcF1M4th0YBV0Qp7nUOax7w3Cnfp1sBZn8trnO2q+wUS1viIzlMFIZT4MplCbj7XaCHc
8P/DHb8/9zC1BAZgGu17SQYNNoop4mjlPNWa0R2uda7pESpzZItiZ4N4jcinyjLepHo9ytmM2gjN
TPUsvd8a/yV7ER/98H5crCfmGdanI27PHINlt/6LoGdoHmc6P38lLRtSLFrBuGZyZ4A+8iH6EIgJ
VgzZjKRIC7fkN32DuFlx14rYWTS69cngkybjhp58TzrkJ0jX/doMhdBOKPYgo7smSVCCRV010mTp
HBMY7qMhtXJ2GI/1S12flhyxCqO0NcPVHgAvnQSQouUjNxuV4zqDIGBrGrk4PKC2HLC6upDECuFx
hkNph913PhRekjqrs3VRy8qiL9WPLXPXnCA/WZ6J00ulguyKbqrU1PDBvA9f8zLPaFICw/x87G3U
a0Es/2Gnffe26gBLSncB5QrYlMuLVPAnE+La5Zeez6XGrBUbZufQpzAXB4RH/zBPvp8cKWG+OTcO
HXO602+ltc0zfEpOwosArvgi8CDy2mYeDglFPcK7U5TU9m4rzXXPnDKZLXHizJnDm4mQLsZShoud
p9oC369odXrk6f281mccKUP5n3aZ0xha/23FEWI1i/nt9io703dzWlE5zg7WMdf3ulJhR7ytu2B1
Tk6AupYJQsFWzba2Zo1pZAUNQ1cLo4txWai9YSE1QUo1mbwjoSDIiuOc7xlaQ7ZBXoOI1suQ4GH9
a30SF2w9J1ABwnjewww9Qf5802av3Mzy22nomtqUfSPeApPjD/oBR2vnWilF8fahMUXkBy8iEuMb
v3eohzIVmQBE4i3yt7kgS5hWggPvyTWYJ0U///K2oWDtNnGtn0FtyrqUPMQa2FuzMkZExO9hdkHW
o9U9QMxIFnwn6tCFafnBVAIn5tJip42zBOb1OYfDOVkNJRRxSrNJAni5MxCcptk6mrTLW2L6Z2Vv
pkwlpqbZl+vzkvjO9pWpei4mAmzjjlNU2E4iKDzV4vkbI6PBLcF6l0JRvEjDBESYTm+U/ryoZtQr
P0Xt1R4lwNcFiog3f120G0Gyixawwm1UZe5rxfu/h9zMWLaOhgVZAf5fGBGfKBTapvd4/QQ3nF1w
n9GIYG0BOB9s3USXwUbYA0OdhLNbO2gHiAVWFQfUzZq4SSaZq1aDS8fkzp7o0jbjdQJ6qauzB0LB
Wt+XzuvN6/mhwjf8VMfPH2F6bGGHi+68t9Enwx0uhHSunIh7bFu/ZfCIyXgCeCiDyWiy20Q1WDCt
uswUfaG/EEDkrs1Qcc4/XWEM33XDMhvuwailsBjyyWoYmXvCrD43547RnJRIDL3u5QDHYL7/8mOc
Yqd5UGOw5IT/RBIsDPZ9ya921Xzy8D7Piv05O0vWe8XRCJ7yiwzKjVYCpn/3fMKxo+3z3vjpZOAl
ydOGmNPoqB136IZnTF1ZS30kw+1Z+29NvYviZd6ZxF5VsJPutmziZKjlYCQA4L8jQUiVBL7gf3uT
Jsh51iGL6Vt+9Qy/cAOejMh3DtvNlqIE5ieHHbsdUjR/OSVfPSn3IMJwwq37HWpwxse2/UOJeYzt
D97HkgrRcrhV3k2g8w29N1kqikRooWZkvLtlbzY12rgsYvHYOO5myt9TuhnJILt5fnfMHgoP3xqg
mqQg02/pNI6FzzoyQWzxFgtC/VzNcI6RxaxW7jfmZB/rJV0GjUAt5Y92lhvFMQ8twT4l1d1/w1sF
DGjiKf0K30KvUtS/LPUZ/318n/Dp0iSYlxMEkj/5DFqUhkdsTCeG97MkjwFjh8SMK5wAVPLXZNK7
j7zP7dEb7McR/x4GSlALXEv8FrpJLZWe1fKUuB1rULY2Hb+pUI+RKurn4DhHM/w/dUtmYgmgOy7G
pB8pdJxg8X4JZmvBtBxFwMr0VHjn1pseyC6t1O9NbWzoTEWxlT2bPIg2wezwhp3irP8iZhHai3Qa
Ev8MvA7m0+lF3jdKZ1XGrfjf+EXrYFfT8SQYV1F6AwIPaDsnZf11XlOc0/x+AHfc9d1RstA8pADL
K4XKD2Px29x26pXBhJOu47PYZBMCGba8nTndf7HsF84xmZK7HYa8z59rkVZoZdu+EIIVO42Zrb1V
Z2+TGuDSW0nAAUwmo4nw6GbYHCISmKomJltpj1sgE6pW+bPSzwQB5uRWOZzpHPQ+GeJvjA8FPzo6
VAZJ8FvJrV1IcmahF0HcSOd0K7k78Gsss+g7tJtREIdQeeHf8QyU3aGNPhvC1wp98FeIwzZ4TI2/
VbtxwpqvRTt79s0ZlUFCmf0EOGqZi5WljdZxFfi4TZLKmGiaHyUC+qCbRPBhN+rrqMcfBkcc+48f
8ktqpB0s0SflEKcE91gqQeVpc1ktcXaiUTmM3Up/SpgRsXiAL9XraL45oFsDn27eFSJG2jwgTW83
tmLFrvAVlOr5vl3cJ6dSB4Xm3L3J9/1fwvmNKu96Yxpabge4TzU0R4YTzkS3CEwsni9ve0SLaags
lMjVXjQCwcke63w9s6ao9TfLOe3Mnxxgj26on+OTDERffZGHPChrC5+hvW2NV05jFkQd7irsBIjZ
8zXCZM8u3w4H7rlxFSOWQFafPRcVQOIGk8Dlrdo5rvwhLls1f+NgCXC6opfPkMDQ1bQO7P5Cdrn2
X0Rpxd/X5k9rfUTAuoHQmHUgB3u/1kgomMllQsjS3qrKXb/bhTlzEWi64zOzlHtVQtRMUbjVLbNn
gbFVHELugZITp1SHwQWX6OMYWCp6s40Q/uIiiEKrG6EzHGX3Jk3E57gRlpR5wdQMWkhh9B6TF4Gf
S1y+qniGkNWxkhL5Jv4/Oa8cayiXVsfnsqghhTYsSTfaYfWtiDzrJXlU4eDneZrGPWQ9Rz/p4J+y
Xc9CraLtVPMtwQShBDsmdmjnhYR1I8sT8G8htQc0RA2E/eRSZonqQUiY58f+yFdXaV/GcYyVBxAY
M7sDdeo+eVyW0BXyN9hMIRkNSKs1/3QJo9ISiH6V5pBvr0a+TZ89hJL4VFQlccqdgp9Q+E7GeWIA
jyLPtCSIHJJnM4PcGdmSYT4u4XIqWo9pcLYIXgoZnor2JJIJkkOFFKv0rKdghkwy9xRIToVXRe6C
w2ZGPBT38qNLZClbZ9jBk+ckKEPgx6K7g1UXBIIAVlW4B+k/M71d/jBGNBvrr6nbwmsqgAoJlQIt
v9QWo1leO0Fj9/f19rV7oOhpEJZZkL+WJubNNzTmES5kasNYhSep2Vfndf7Xaq0B5nJE62/oUMIa
Uw7xFSsMlP90JHjgR0T2KmjS8p1VKQakndFkac+aily8faSg05K9xw9RrzTDMZiudeFhhEFR5di+
KinymuYx8h60cjOSdV9cAci5vg6I6z1wkAzJyhjBxRnQj3DTtwUf9ja89lPFIuo1ZwItPhWCdqhw
GKuAcihLjOQEJ7go2pPIryB7FhRfjL6LjQxfP3jqxSoq5iMhxn+Mpj+4dDWr9JWg6BBtlVGMR/3U
axncJSUYPg/fmnnaz26gLeu7S2BCMXYdNM3B7eWm7ug4rxv0pgoPE4aFKmDfNZdU/lawO8pXSFmC
hejr3HYQbDFphVZRDTOJnNIxUgIRXa2LhZh1UOaVZ3gJTfv92kn9RB3Fn3+86NXV3gQFIRWwKcdT
gQaHqJqvfj8KCome05zEEaqxx9PxUD1SPcmGsjnIp1oAwkS5Qqrr60DEPde105/2YfiuTVMXNWyO
bGCRvrrWiYBbMjQvkmKo1weplEwZJtvgD6u+PKFVTi2Gs05zo0t6bxB1Iuo8/S/6QeCBqtHlBsRk
lJ6sbTbXmIw6qjpyt0g6L6Ofub0rHRcvPsy9h9bQ5Q+G3PYTdwuamJgDkKROzD2gmknpBGUtPrWy
Wca05/gIEwmyd820opmxeIjUi7o0kvAS16ul75uua3qXpOD07ofXWTm+Bo7KslD2kf3dnAYhUPEU
mmEk787LrJ/MwkMloBWwZlG+cVKj8rt1lFn0dGlQxqduqGgXegjJVkRIltTGmDV5sGehiFgadoS7
+uroYsX9lUEKppOJq1uo2oPOeRbMo/E8AdTMG9zKzRQVpHQ4hA55JrnCOAnv4vIRz2fn+Q/uRdyu
Gs/Bo1giJJMFrkCPljSHlSYlpCzfr+UZfMcBoaeB081OrXce0fJvKSl23baxBBMdfhBAatRh2LVc
SrD3CZWIzV+YNgkv3g2lBKF/b2I1M7Wv97JvAgv7oXZU/BU2lqUuSEdQY03TKztm3q8e/59ISK07
q2QHQrO5vT59QXh4acGkLDPueolN2r3jUNw80wy8s9tH+S1GtU/ISPfk/q02kFkYE25FXJJCSuL6
mtiPaWt5HreGfqwKxhPv4L9tWzCm2OmXkdyrxlVlDjdcWKslciRFFIxjd7MoCHwB3v1eEjhFyODU
G9jy99lSkXTcAdfyIP5nrn986D2GnS0uegc/ukuiBcEndVnOw/Ri9vEdsAefbx2y2CVMNGVsdMgw
+mszv0cNknO5dbEfVMPrRdIBFQZLeXPm//fe25Om8mBkhRJvgEjbBge1vH1fHcrnMovDdDGhlPHi
oc7JnIVV0UbnPumU/+KmZ7sf2HLjW0byfV5QoK7ssKgUlaK5YlOCwRzeP+M8JTA4Cgp0ifcajUG1
nINNK0VGTAQczTrcuK2toOYCrq543aO14GQWFoUaE7HjKBHh4E7jm0P0M9PEaWCfbpuHjnbYbMXG
xN6seVVC6S1g3Ij04BfrebTSRhdqhvJocHk9tW5c30P5+kFhdMAf8tC0Pu+6jFuuVxuE6vBth9Vy
Jezg7EA7Y9mzzHA5fbeEkj01u7i6/ZTfek2Oj9OZetuYxYlF46k/MFf8SA1hu+FYGeZgpkhucrzM
W8cbbWD8UCW83He+cihHh2wfomjjn61KMZghSnP8qGpR1z+Y4Lvzfcu/wb2XFQ0LDXeVwGTa8Hmx
BkwtWADbKz/SOvGbMi6SsfWOUHh1uPs3kI7qwM9IFObN3v9cQnVlx21MHVJ79HSuIKkHgQH7xPkS
walrR8OGUNmguASXDcjCTbCEv/kGfIK+n593qjuhQguYJm0+H3L75rVWpVA7trGr3ZCsRWmq5l68
Ouvm19yY5u+DtdPv8xrUr3KMGfFX5pmauib6xJTeb8vsMkYe/eQI2VQ6EHEa7cm9XBlATUA5pbk9
t+UIqtxYtvo2NukFa6TAvQu1hevknfw8OeawEqUYQ7nDdg2X4/XBmVB3AxGhNbx/xW+Am3psNSaC
uOD8guwV9n7TrM5swbXwP/V5b2MLtLdcRblPKyJiCciwJ+EImsaD/bcfzeaIUowx+mDDcyogsnEt
ALMJXxUfo0dXwQoUKEcaoh3EXJPomekaNy26qkBgt8Eyg3ri74HzIDVLhZm13jFExLG01IroYmv3
/r5ijb0J1WVSq4SXzv7yeJPNNeAyBe628bshZLauquNmQzXfxF8P5TwlumM+thRMxLjvnZq+rPIH
GEiLrw1uZ6Bx2rZOIfD/ALJBD22GoaE4PpfjK3xMFfDX3319wwEeSSRCAK/+jGk1FlJfV/TnEfli
njmVEXvyGmS59Q+BXh5KugOm8fXCxkSjvbS8qgvmANAw/6KlFlBtzUQJFRfvL6E/fp1Pjt7ocn8U
c2Sd+aVv/hQ2LQpnghq8zqR6EhperLBLjVFf207aGRMK6Wgs3sJYAm76U05eoRCLlpOpks4NyyRH
khsuG8KkWhk1LDWKNrQWUdLhSj2d9pwNKGBaNAV8KUrMKVbdGcvQdfCV2FvY/UmSJFCpyHjoikzL
d1hpsIsUoLEFZSKidPP0CfdkT56dfGerRR5NNL76ISaEfJ78elwYsVEhHoejuRAqRTCL0u6W65Vi
B6J3iMxEckv8ewpW8pnaE3uu8ccfJB7klL65BZfoz/wOGErhlnIhb+bna7x7uK/5HARxsC5Urut0
cHMRM+BQJmBX9kO2LLPD9agAiMPenfYN5blZOlfM7j4lsh0mrOOfAZIW4PN27B+/q7U26+leXltw
aVa5OPr39wm7oAWdOsn3KvVJyEFMnDQwVoLA6aYPXbpl7qyAuHsWyRG1g+FjAPSUwvzY6RYS3TmN
uQIAGLKtZG5pFrJyTwEAeH2rGKGjFFCR5RYyX4N5miWXlqNLBPAFRl8pxSVJsS+efXyzrVCwoKCb
rLop8v5L9FdNKJiF97icawHnLYVchs0SliWJcNmkGHi/j5OwnayscBJLuejp+ffVAWHK987q8+2m
TjMEOZ9wVLBLsC3i275lnxgi6cFhpfQbOFrTaBav/ec3Li4F1RirfGIsnj1m4HdjxeOfdfkXE7md
x8/iuownylR5k5K5Vo4HccmI7AoUToGhvWeDiSl48iJ8ED1tjPaOVc9j03RTy5pbq12JOzSyzLOa
43vBGEtKu0XmRQ7oMIcAurHPhdNsupEvRO35LaoNviNGLcoEru+d2aQYYpvAKZCoR967/YTb3Fn+
WqjN3yXoWoBQzLfwjko8hqXPXoOPMjJB1oGjCYyHVdXejO5xKxXCdhQ59zfPSrqF0yry06cmohnh
qsF+w6kxo0odCqWCI3NqFG4wC2Olph3bjoD5iedww3W3//WfqFJF6PAwhpFd49Gy76ZiH1O1sc8s
PpruWFZ8tjs6JISRCn8w6dWRNgbocMTEKbKoXVJrpOwv4ECRP0Vk55jJVAiA3HCv6KRX0Z7cZS/h
hB6R3i6YaEPcInkwwBStEwlbOxxjTVX0rjgZCOpM3ccy1bUy9FRwAo3JH4Y1MhHV9NGQtac8uaIu
1wB71wAawDzRYvSFuKn+o4VPOVpcX9u2gZ/ePfymN/7q0f42h5pJuHtchpWefYKDqkH4SqdXxYlx
hiPxpnKaXbk1p4jiaWJ+VLggSBDPdWk7UfrbFJWNFN7OUY0gcbeWOm+OYDngbH7z5fTgGUHRiky7
zfHxsrjkNhM8tM7ARa2osZ6RMlDnAuBzIltebXelG6HdcGn0mv5txUefvo92O7HkGo/Xs7BCvlrO
+xp4kqQ/D/pGKN/IfUPd5+mh+uCC1VGxgA/DzisWwiugiY2PRrI84TkmaGfXj0vCwCQGUodNDQ+9
GWMsWqBg7bka6+pI5It0ROmxsdILT4v1Noa0BLuChSIcqyJMZmf9f/SaHyPypsC5cvi9EPOCNmqR
0+o04bVWpMaGvzT8c8hcvFGRzXTEGLKPKTFLuSOPlHgZZEtRq+3spCyNTEAkL6pBKWTqNGI5b2Vx
oUcNSP9DzCDb4jVxqrnnvbXdPvdvuV59NR7Gd7+KiF9XfGK+rQzHanjOSmt0GIeZa0AS2qq2qIpq
QqUq8mPMa4aZ3xjDn3qtg1mkEkCUhJr4JPBPM1ULtBCvdbG5TywxvREu89oqNecMnDGnGG+Tk/Ob
/tH/jbDleKjwS857c1JnlqCsHrC8mfaBNO1WjWSzEBl10X6aEwaQ66XazxjC367nHoGEDf093KmA
ZDrANwTiwLpxF5ynPKf1NKsKOVtT5NaV6ioDtpIrkSdaVvA1i1IuuksL7cJjqvFUVb8n8jPRBIo1
TRtV0P4iXTTyulODC7ITiHQdknHlxhur0PtQt1rHILL2M9IXkXSmD+3h/vdDgFkyM3I3AFdLhmB5
rdIK0p2Q4NRk2TBu8T90grE43A74Ew0EKKGbOX8VWR0/MkAzKFddaYDZRRoCUw8bTRHdV6zhOVb9
DOsi+36/n05F+AiYyBxgg4yL5PUxETUexH4teTq9flptWlpyyU7++ulywTG3OvbkGWwBvzYfCG44
V1Xbdj9ZKE2BVS9zmJ8QvSJ7YymgbU7mG7OR6JYcdvo7fp+2Jz7UqCUTAD8HL4TVy5if2CSp767a
D6N2VoWCmXwKtowOQcU/eHGvGAyX7YMXGgJMSjLe9k/mHuNMlhrNF9cLUMs+ZJ9PpB/7q/xLiuaE
f+goma5XptW8N/Uyq1EJS/Wh12vqOGTt9n8lu7PXfK/TDjpX1mRCDV7ZCPz4/ot+DQeSj0prcGEC
chQBn9uE4KafWbLCvZh6ce8jD9NmqdT5JCYFZMPGvmYbl+5nl/KqM/7SJp2RYi3oeEm5LHEyrM23
Rnl0O9/hS91MJUxDrOT+rsYm17ji6JoOs/hqBmC4IivKLP+AZngXcQR70XREA9Hvxr9iVDTPuxkL
cgOnaO1cxQsFMUWw4tP0lvwrzgxw0tqUcMUY3iNs8CCIimMPUkRAdnepTjD2Lmh+UvNwY5Cq51jX
lUWN6BHksd+NLgMJUROnuS4djvH2v8JAYapSetvQLpL3o76WHRArr70jyqOGBFe5cdIODm22abVJ
CyiMTrVxfuoqLeEognl7JwemOdGBgLpn/tb4KNQ40bA9P6e3m3nM8Ht+waBw24/1J4wwzTeWhZ9I
n/1OMF/8bdVeseJhzVqxgLM1i5o1bCOKL4VIADNUpoR8DXA+1BBfgMcUck9Yrl/BW1B0cLVFgbiB
YihSdgK6+nHUndPTZQiSrs/xqIvtROxJx0r/XApWLtTOythaeiMFuPay+t5Kj/GVpiSCPLi5ISbA
NQqIMwoVbq6S4hJefGODB9dU5tCvszprAhaRZ2FKyfLCZ3kfrLPn3qneBAB6Ol8hLSEdiXS3iUbY
ba860MbYTqwItE3jO8ieQJlOLCtXYCmK7yJIP3N5zzcEVkEQL1nqRhRbHEqGcdf95hkFTuiIxMGA
Iq2Qd055D5BT+xwim5lj84mBrdt0D9OP/AtVweD1UCe8FZ7AuiGmMiPWp7jWvoiB7Hqb+39e9Zuh
9q78JZ04fosACA2srt8GnV59TLBsTaXs35cbI5aPgPu0Hh3BydTRhj+An6PxT1qa5fvbbexXhWeS
BJFfsnRkWIT6l+ZFNxf8UM5wd2MoD8+Q+3apDp16fGNK+Hvih/dfJWGw5re6567v6gXKS9aXsj7T
cU/vME+si7p8StkO1HzKe5H+2ROQG6kjMw7EbZMTcdkLjN8BjGyxxiyRv0PfpeCghGwU0pszUhBe
pvfv4AHvxPOyNa3GLK4/lpAQG2NXTM7unL7E89ZNo8G3zvtqjmQIXOQkvNOw+CqYm6MgGsTzVfuQ
hwDYpZbxlAEnHjtqUXrPVuBXwtcFM7AlBXpkZtokndm3SXqYIuCqbx5PzT30LUTGiToLCqxN+XF8
q5j+YgfU7HS2IyS/taTRF2L+nqQkUV/8+piYopfAsYdR2Yshyx71K4aTUJzEWcwDIKTe7lH/q3yQ
wstVQdrG7qWRG65GhDhCLkGyKUHELafIO2awgHEqGaazqRtWYqZcC4MoB+aoHYUFdc2hq4nf70yp
GVbfT4Z+hBdOycCmwnVWh6mBAz4AL9rybh96Y9EvmnHx+4y7DPVD5+N22OgKMg6DDx1+cjunaLHq
7TvUjtCGXl//vSLVe2EYeKrT0KRLvduZLi3dYGhl3hm/sVDKSngpaYQwhsRi8PY43wO0JbSpQbDg
XnzNkpxtoGe7L47/G+Rl0RLfpcvLAk+S30HvXbGDPbwjjJ2xzmuWNuARXylto/hJlfgyyEbHrJbp
qX+O4DLw7kIiNA5rBjNoJrpmBTuVsfhj+fdjGFfNIVWPQm0YmE6liehAt4m19CaWvYV4Yv7GD0I3
xJukZHuELTkHQ5Tk/+P5NJvaHNWhzObGSrNsebA0Wh7CqX+LjDrKgBhnBC/n/ULOICsD567ZP2ee
AP49DZB2Qjb5x8ihOot3N8Y5QFG9DkbUDHjoXM2ZITMYsemIRThc3+6smAPNr++zmhoFbX69GXuD
FYK9/4EQucH82p8HOcufde1iaKHTw96Un0U0Cd9gd9Wjgap8DHd+GdCK17NniRlloj0Hq3IXqd8t
5OktN07gAVPp1HyQMSd15gdeDlYQnEFAxVKvu1pk2ChnOq54YGF2HHLELirUoQ2oy3GdbM1LHbLe
UjMRYA2NX/SO7o7c5NgLp0ym0quRk+IsdtSDIaJ4Pu+8Uq/ERPMln+kWNjN2pUcEPgNAqREYmH0L
U5FIG5AanSKDH6dsE34wDT028m8XPRemTSF74iGDYAgHBNoQw/WG9MHzmGKjJeY8op019C5ajzHV
5aYdi+XfheRdLqiqQzwTAiV1pycpF3GU34bk/RohTtRV6R40fhz2L6Xpf65KEg/hURcVPZHC7uPQ
/A92goUn4+1Z5xBy6r9lZ1tQX4iAeiK35edyyICyYj5z5nxv3SZbYtNq2o3uzKkmtJRq7pfNdRZ3
hL3DtkMWHaunppoIhaf6KZif96eD76lZuERzJXXReZl5wWAYhKaoHEVrbCwnyQxcEhMU/VZvO+Qz
d8Txg8K3J6JMYE8zkxsMs6hubQvyapaNQu4RsqzswNRvGmw+ssRpVof5B8Q7sgS+XQEwud58bMJl
5ApoDnfyHUudq8aaFqOleiZ0XlE57E3KXA3wOpUekwUxnICXLK4G4aR4honqBNXayRDRWNet2mJw
7HOSzq+1PArTCSOc621Wo0kq0dfXnenWEtiyuCdCGUsrOqsnoojdrrIKc6m3yBdIGVMfmA8njA91
Oz5KzXa9t7vwEm/GH/2udRdCUEYf013HS3M/5JdXky77tyjiWGgdHJXMVZlBoTa0+a3MrQ8CT374
DJFc14mf5CUDPeNRWHdZCO4vgncU2FDRbsbsI/BWiyGzBBKH8lKEWEjwuBynKTNGXjIBLlTob1Vk
+Wx5hoMdLND2GTeDn3q0GyZOrqfeDXQMG8htsW/Ik1blf1o0aoZ7pg9x8LYJKPAfPpUAG6diB9vw
rOq4z9ABXB+WOtd0MpNyLQl+rtTQeMSjl7i72Jl1EvlefT2J964O+nAkh2kfoCD/KFV/qjgymWYU
MhusqlJb9pZm3iKQxsPwg3astyVi8QdeR8gXaBerC4qN5VZvjfxeC+kZlbqFjIyU9NiCkfUGQPEF
UyuOfg0hsOArTLbODjT+jHPYIkaI2OvmohWNTjLEAVqZn4ugS6TOKjq9BS77KPccqiEkZf6xX2Nm
AFJXimYkaTHMA0B/qNkcqFYq1Xw20MPn+g7JCEzruOfgHkElL3nBIuQXjbZt9sNoJA38/fe+j3Uc
uUiTi0ZiNe2nkQ8SCKF48QGa845MqxYgwDRipn35YEtx2eKv3Mm+Rj8arEvGsGAArAcMPUjLvyBH
TZW8N8CdVeGuosDxcGaZY2sSW68HwSTEAfgnzb4DW0Hty0xo5mCqlUw8hluxv6elUKFLgJwXyfEl
lTNGXGHP6GnQ0UEmQhE8ooXTIe2rqGL08h5VRpOwU5ODgtI0v6BGWo0BUQRSDikqPgjFEj9hWfBY
OFhhty0Y+LC+z0u4UC1aI/ZX29gzlEmy91S52V84j8lswg9WtUvaqgTYwNkicU7fSzbqXogGQnJc
mT0M9TYUFDHMJ5wxzXP6bOBgMsvhe29fJT9kUmrFklpDeraxk7LffjoKH04l5KV1/Jnz/+tXXD4C
HGuGlZQYqzW7/XyXRf4dJ+umH6tJQjVcCTkVXRUoYhiTtwVvrOhfb0OlMdFCm7hSOJccdWrQYhxb
Bi479/5vF5mWfYsjFKYKGOANCc67Ojq6udef4BQwh7ItcsEEkehSwjyPms4FINvoapX73t747dVZ
Z+iXvZFjfvJprUty/Lo0NCttcYnAJ793x72VL+z1SPy+z2Yf+SAkSHweOVNivFzWnWmFI9auXlOs
MbSGyIfCGIaYu40sLOfIOP4oS8ToItjtAdsd+GwnXO9+O0UNfKDjebthbN1yVuOf6uiUi6Owho2d
mTjpU/c9uU647kMBldYdwkA3ggvjMenpjZMtXyjDqFEh7mKawrKPKjdsnoXtzBhLNfNUtsANx7mR
kX1Ey9k0ZQRI66NbJkb+9OsKYxNbd7C+REWf6OTuGYgVu1/wzYRm39kGUGLH/DQphgNoY/PNlFyf
wCaOzUIpE/WJ98kNWY89iu+5XlyO7/0pyhc/N37q2VTeNBJaMrFCoNCz0Bitgm/NkSYBgY6xmyCa
K7ryJBKAWG6CInHEm9D8hfaxF6eWiSfi/jpVuuSLghpe3M2AGLUvEUOjWsc/nc+BQLo6MxX6Hel+
fTrjvqLEDonoh6tg2VU0E3++MgbtNrknc7GWbKJFnFQxlijKjeFGIJZ8MReJCSPbuEzIonpTc2QV
bUcclwh7NqsWLUdkiX9/Chhqz+rFASF0Gag2jnEdqRgjaRUow6MDXBHu97OZUK4GYXOLgUxCbTbc
9TLwyzqKhwuNFHzeLfcgUVX3CipCwn3UWU4CJgpTN38wXxI3wzQ8cqsMetHFh3hwrzCA5ztv83mm
CmSVKHFSUe/lizvVLtY+LrzFhAFu/Lfp/LVDr0oeOSvATKghaB5YhQ3vrYGRYFVGwS9kRIZ9c0N9
Dxv47niyq79z63RZldq34DQ58dbu6PPA9qUtcmwPy9NvJCslv+OE6gEu7eog0wnuwZSCF3T2XEuv
FgyDOdfxBdF2MadtrbF4XGBYmWidEGUa/LLnqJwZe/xmW0MT+yGhTk73STu0hr4EhMrJ9LqQQZ5g
do8YJ5Equi24GJUoGC+PekpjCw3DAuqd4XhkThvkhwoXAX8eOP5ybTQlU7lLa9t8ct87laxkgQMp
Bopg7kIBPV76nggKwrcCWCUjbh4Uvf3N7mrRFMjimi2hVPdjPDBXBdevdm7NJV/IMA/N1DlpdrIH
8C7R6ocRez9yRjmR5Nj2V80OuzLXMKFuWfZUMvsur1We5w8mbKUAs5IpGDbeSFw0+mPX9gsUZC2K
nQaZkoIIgMz+ZxatwS6CTF+vpnfuC4bI8bUM/uju9zsjvO9tWRxQBMvzlrYXrFQxumnSwMEuSM54
HTLYQjpdUP2SnsShZFVeBKuIx2eCGt45K2/P5CIDIbuDI+bxMlDxxtQwpEKoBvhOQ/rP0lsdTfu/
aFxueN1rZjU23e8els7c1RBJLdNmGb47NS3cAVPikCKObUeHe/NF2uL6CoYklEKVxnexUueZEhhR
/Vn9CrJLv461uJHngF+Bh9wMlpCEeK0e/ytj9njWoiRMKz0Tk+KVC8iNyxHebOzPo5nwtWwQx+XM
apizbEiq3u4AcAMPgf96vAJpSFOt2csrnmmQ8MPWezWLHbFuGF2kp7AUZYRTXIkdz/lTAnVxF/4H
udxMhOfW2cy6EwPWTd0mfrJjQ1EwRE2YyvDRK2Sipw3pkpRrDf7fHiUetFs4Er1sZw9r7eAemy0N
BBYBGJ+l13PuM9j1rQafuBhmjeXvGmt5D0N2+NU/qe8NyS2xIcXjGn7Tm3zFRWllLKFTzo3X7MO9
QyDvo0xMN7VcATqHREIwRheWfSCC2ct+qmOwb1UrxPzQC0l775OWJRI4/WYgUHLa03u09dIkEavG
y2smdx8bQ7zQkQCMeFo65X3kKAi5L3AnnX6QGnckyN+Scu+Lh+mYp7qlBTsoLFfrknHJ67clxj36
4cWhTX2Poo8cHKhMhcMhye4ge5md/PJD6vgV8CS5vczi03q9RHOmCGjh2Yn9SNba633wJ8RM2+eu
I6erPsTQl46EdL/TBsNS96EtNUtPq4N8K2wPalMgnqb+39xB1s+yYTZGALTgDqSXFg8jGikLJ7EG
IZMH+rizmynyQEazkOBH1UsXfyEbdjAo7malrjCGbLwUzUouw67fxoQ9e1yX3Zrnzn68G3i6bEM4
d+j5tZOmg5LuZJyv/WqjvjreP/1+v/SZ6qBuj9KGOynCSpShpd//TdnyHZ6hEozO8cwoYLRZjbI7
xu3Ywwlpa5iMQ3Pd87ZqUaVHEjJlf72WdBEqE6ZMnicpI1xwV6FhAHNhJ4eVvH+9C/+rFsku7oCY
Pu1wqMpbjUD+g+37nYFSdEfEQHd73ZSyZLbGnQWjipFM5KxEfkANpo4RNEwPl4wk+lhAIxg+4xU+
eyLxHU2sAnDS70V1w1FHy50nuxuAmm1PWJCxdsFiAHJfgFrY1ZZGGiIGwbpYvPQQuCirmxpR4qi+
+ebiHv3DVOK4gqmlqI6Pq3Y+CM17HEd1OB76vE4HPhvKUJ7XckvQ6RX3k++/iVJembZFRdJI3rCq
ggcIFV9cX/Tk68m7vGoXXgRl5SWmfW0aIR5YavK1tOSkzHjdkjYZAcxJdLc5bqV2lSA7uz2itjm2
u9oOImG4S6smDvULPrKzY5DafzcF3uz1zv2xfTLrrSsXge9VytgwOxO+6LRJFSWYILfcFArgVG5j
J0tC+TV7hwVcGU6OfCiQrkZmBE2bkaPmQYtCqevrGKP6KguearN2GHHjVW+wDmAWRu9Uo9e+obXQ
g1IwmrucolLruX/RTBlXFq4EkSYHxjFRXTyQNgGqUSqZiwpa3wShzPtp2MZNyIkrkBlvw6m+E65N
Q16Qdd4rW73Pu1CYEff7HjS+KdbWa9IcW5j6ZYzFvp4tGpUGE2xIPyKhA28CyHtqYd02zamjiLQS
IDkvKxRMWCHaO6ZeG7WyNh2ju8dP5EW5vpvndVzYjFXlEaabZ4s5BOw3+y9a+QWvXgfM6rQfWii1
u+v3RQgk3Rbt9ntRYICKVigZFkTkhqfAETVz8aHX68XrEWkZ3m3VjfiJtT4vBbkoI0vrwR/hrg0W
5xKjrme8YBZTL+wQGPSbiAssrctGUXTrOmC0Lv5dyaUVX8rWvlKj4/KAjZgM7GXxTTGGt5PJ0UeN
fTYHEFWbEK57tilJg1M9Nxvo1DHzX3fV5TPQjnntWFQaJ0k+vZvML+mGFeIcNV2BcWH072ZfsboF
wB+IlaC6HypgJApDZJ/hp7oZf5xTDFTgXRWwEN9vySJMnkFpK3rg4e/z75BxE27UyEtNiQveP3ct
JQ5WS0eiq3S77FI3I64kK3Jzf8219UfbjKg/s0046pR+IyP0AustfLsbp0MSTF2zKW9yryuIdIoB
4TYxiscjghpgjW5uCIiu5ArKWjGU7Jph5YhE1/qD3ak941USHtzmJJ822qPmP96pC3hVCx4vvctJ
z9HW4ncuIxv7i5W3MK9Jrc0abRgZgG6TF3N/G1LJKMMe9rs8OyReUdJPQxkaZo095mJLP7JvuSVL
fVHB7aiEOPpLTSuYDAsPaIWr9Jx4ABy9SFrLTGhdmQjLdgGK/VGo2c3Q+sRnP+sBodxCOcu4XBay
/tSy8PMiQ2ymnWYP/DsgiSHAQ6siKvEIboU1UYgBn3EDke1do/yWpcxfTFzvbYiWIV+vp7cFnxXS
v3Ky1ehhZiiUHypdpFezgeEfmd/FNSnjcDKwxxkeWwSdAjQ5/NPzQAmXdVpYhpsPQLFylfYdkpPU
NJ3kjaCw5a82aghyV+CS7xLU0GJQNN/ZrDgwZdrcQ/JTyM62rjYK4F8gMAOXaGPqQgWBwAgxzv9B
VzBiQdoxyyUJM3mKIJXDAIFb0AcR4cGn8iVE49yMpbTFHoAivJYRNgU3WCx75WwIGe4AdGWYkU6x
37MBBbpeTvJx7kZ824y1y5fTnJliDTdQx6xxNe3NjDsj/vAUOQjE7onB4X3CV0uhtn8QLGSr4ffL
MIBbVQEIFGMY3Lgdm26udhe4QpIgep5r5OplrH6uRtaQbfOLGf0Vi8fQo8pRT8yn01+Jx+hujKvo
SFoooPi0acCvmor9/gVSsUm14KipHzfWfLIGA+w3HADpAmI7vent9DJacKxu0SN807IdMcbDv7Jq
F3ADvXwRLkfT+MmTwZrX87kPAPEcBI9RSSsRpqPiPDboshrsHZph6T4bSnxF/FweLOs3o40JvN04
CderX+goyJ+Ac5cNz1iK3qVrPlDHDOezyvZuauUgHcYTUhrdFuAISvoA/IFN/z79YNyMEKoRYOWZ
JxEx5WoMuUFNpR+euh9dFXT2ml/6rnryr1z83WqF/I2NY60gKKuYUkrNY6gxrUAroCmRBQavtk6h
pAkU8cHKSK9MOmZH7TCxeI8GV0dJYLc+CVuibYUwRIkat+GLc4bMikvMplbld+/gcr2HTFNWcjcp
E/823OntB1ZlvfZ6qLwbnCR98ch3C8F4uBTkBZkTMrkcLAd7naFhu8zzJIdDOdTkrLXVIyr5cmM1
erzfqzNxs8HcvUxxBX4SzL1GW1b/h8ylqXtdxbuvRq7Ip52yvstR/DqBOZBWF7nStB5dvjKDSyHu
roS3lJZx3xpPilD9x9PCFQDmwPk8Bx5y8FGxnyP7z5CVMX2Posh2Zr3Dc+QW3OKATnEot5Lws2nU
HZIAGPL2LE4RY2S/jVycd0AkhsfOpnwv9QM9PmFyKAyyhq/CDHcG124NssFKNdc0zmRSNdMhQG+a
0Q13Cy887hmp85IHiFjdEErlejGHg4aO4OLEtnZ3G6p398InqV8+x8RiVTekZ7ZfTTqQDc0Mh1lw
bAroSPiWLiLMWGhaUs1bGc0K3kJ/rQsnILKkLZu4KxDkaXHrmoQhbc08a2MmX97r/KfUFFelo2vp
KvxP2ujy+Ov5LOe2dgqNKihrfbJnR8L/BNUSlhdBF67pe2CESpz/bVKmdI9kXxPyLehiwtYU7kn8
SLTv1oEctqT3dRaN/omnVDRO4SZmVwTXcLUo1KbRBOHi/MXTCPNr/m0oI1m0vbaI+36/CmCWpGLq
0xCRN1+JjJHWPakEaXxOcD48wKDN9dEHhdZy2cChXzb2XP9s1GatcnIU+egEj/B7DV7hOX+b9ZWG
Hai5oEmiuMaCVLMucKssKo9mFioSEiXlXwKB4FyixevWJeHeHa7+wDxDQvG9DtcEWQ5eCvEfgCWl
P51bSG6rp7f0RfEuLInAM7gmggDcY71YtvN/57ueBFXXVmKE1vnPTozqblw9f22iFzHnRq//YzOd
CQZLO6NrsSL4Bkxq8dtq/UwJ5g9MUSjeo+VkdfCB7YlRKTPQAAlmCzxYr2pucY5kOLX4SufAfEAx
DtnfdDybn+wpI3y4KH+NqIkRMj8ZnqupsRqLjhA7IC+xhMKXkq8AR0jn9s5JfhKJbLthxjDDPcaB
kGLEgbAJq5MhNUS2MZi0lPuRGBnUon3bXxCBOloCM2jxLxN1slwT7+vd/JMNQ1H1ODk/st4Vxati
Gk1TvMgOuVeKaTTfOgBO7ydYTOTXlmrpvhN02/YKNx9WHUSeIMY4pZDzlZoxtuMeO0FMBjVI1uzQ
WkU/wzJwTBZiw3UquHl1tL0uH1OezrLhMJz7SMq+c70fZqCiNFSUIzAc6McHhZZhq5Kz8dO90bO1
z0ul28BG4dOrqYAt28cbhTYB70SSP3ghXN9jp5wbVKn6Gn/kXDi4gaAls1rtygVX2+tY3u7TDn9N
LbXg9INhDctU6ZhhIZJgFygY4Yk1iKNUBouGKHTxLsxAY6maHHszEFvZWB7o0WRCXhQfvVR3ksyl
lJiyKs+TU2JeTscOZT9iGbI1ESZh2zPSG3CEdea+k9qPqV5ocVu80tYVZoXSYhrUSDted+T6lAyh
/71Qf9Fi70kvfyZJagdPgXUfzJsqbkJKODjwTz98MDI2oDKAGyFJrjce2DA317xObdcR8psY9SCm
SzNQOcG5yA80URJL09iQ7mNZFxKxb2nwU0z+OkNT7gGUOYCSNQY3r42nzizIUuoWKKhP8si5c+jU
+L+RXL2SgYLrr7ECWHbTvth4mDGVtEL3oUZgr3n2pZ7Shvb9/X7vn/+dkiGpteo/hFiAr2auQY5L
fI6Xn945Ifvf0+VOYTteEPrpWrgZRO4ofO8P1ov5yrgBPvF4aORt4+w/8wp2QKeOqKeXobFnAM9M
kaATASbhmrq+XZY6vLwHFK9XpwFYzFlxwBEJiaH3Gtn7jsV0UjhYyqM66qD+TgXgfajFwSX0HIAM
Y5TbNk01K7QOvylAlgdrRxlJ/nvzVdfoZ1/eDcZ8yCpAxgRmgStrenEbjnzAVnnw3DShcu59rh5w
o8WSVMTH/aYRj0TEX8mrSKb5JLl6l6oQov/QJ8A7CWLm9QKuSOpnLocaZua23tGnlUhCwTy6CKIU
pB2SCQvASDmEmP1/FYsh/z/FaOwqAMtKMB5CRrRCKrbsa3xinYQZRjCQ/znDm4p/sLM32bBECZi1
cMIzyhXZMcZD2ja9WVPOYdvvbIdIHI7k2uwe3+FCNfc3+v3in5bZWh88TQB8kI+40xEaHneRvmZD
Bp8vLKP0e8PAE1AXe28bcUNVtm8HsYv25A4hKHn66xaWtGA2N+mWqVmKmjNrhVrXVSgJM5mM01iK
gtGsCDaiE8mRpMUqWqZK3UeMjpKe8k6LOGE7ryz2ZGr2V5IfaMBicNS5P1xmh2Dg1dtHIQgrgdq3
9pklFOEanu6zrPh0SvSw6kohbT77xNTvt1b3dpmh0rAYL+g2cbmf41QUZCYvx/Px9VT1Mj8//Ph8
28OT2gbnKfncWxeCvzCR1dSxkMkstOvfdYyY3V4p/9GgVvPXKEwLF7iB6Sm17w1yPp+O0DxmR9Bj
hZCfInh3OfoWVutJV0xyMxB7jcvOn3owWnEwOJvjEE57WZcMBagv8cuTBDnBVtDR8OodTjkspmG9
zPqpq3eoh8aOXkrxhQzDd/gA4KRQQz+eWLIu7bZY+fZ3HcLXeGQ1E5Pn0LJVcvIKk+VTV1jKqYVD
tC8GdoJN7ea2svriQGpPbQeaV9w9kF53d8Yq778UHO+LBYDNZqfK9ysHXViE4TwHgoPW4b6kL0Uz
cNDql5ljj/48KNkMtWorxE7A3cz/p6FKvw6P6BadQr6LX5mXGxQhP73Te7Vi6pHuWOsneE4dxg1F
Hh5Ohgjx6k6NTuog3E0qwlbdqdKHrKzflrJTdscQ8HeT5Upiqs9Otyy1ff5T4uDg1bgVjRkBFhVZ
CLg812i1t7xKrq29a/DjXWGmo03/4knhoXUtVRTzIzObHtCEyvt/PgqTYigu5jgY06zOXUCPbOGC
HG0CHpd0SvluePtc3v+rRaryyWImhvZ2dnG2TWhjuP9op4sU9CzlYjzZ6se05cSij0Y8SJxIvxqD
vaPXRYq5jcVfmszaPTV3D6HvNhg70O9Lu29jWrymIQs9v2V8P2Zjis10zcFOeGZ23q0SpPCLVahg
2eh7vV08+/dj4+VWQJn5kn6LUkrJXmHXQ3yJjgJ1UpfAIU02nCvfbP7pf22Ap0lQ7LeiPwtIFde+
l6CT09/3rOmn+VMbui4x5Dssm5Xx7CPfnmjUmEoZmua9qHv8JuScs9Qhb7Th6hKl7d/dT3k4bWx2
xWytPL2UoswoWe11Vur0NYBVzYTwWX1i39HfnvGyYqAUZYafNBfTcwZUdt0xDEDRaI4oFLfWVS45
+humJpWDuTvXrsWMXP73EY+oS9ZF+STcDRpy0gJ7s0mLMjytjZbMswtrIxa1KUZhBr3ZfTH/T0GT
qfqg/RcWGgdSIcupj/Z1xnK+TWpRjInHMRBQI0A9eT3isCRx948FoBqNtIQlznNREmZtqz/CEkuH
FzlOODWCaBrHVb6hipjyz83iZIj+kOodG+P9XFhXlb/SNwWHD7HpGN6Unq+rM987vwTM2l7gyxwS
WZto4pM/90jJI6goUzc+O78TYdiyYt2TdvPz/ytIqY71Yl/LzOgqqOsT0b2mcD7AoItSt3RK++Sb
5uPc0xc0ggArrjqLdzlwiADF0Wim6tQb32lvp4lAP2wj6Mdpt+d3Qw6B7nvi6G45TY7Q0hCyre61
9dc9cIhD9S/fQBcrEgi5l2A1xhsM+wa1EioVelIvc1lTk+ngzTTN1GagahVPS1zh2ZQEMDuQOEKG
TyywvtQLxFy7XgM0kX7Dca5Jddebz3jhMOsMiwXjquh7CY7l2yJJFh7STgpvLfc9pO2JNKwRTNxr
5EyUITkFAdzgr5FZTj1aedvrzBKvBJJB580QYosUhNyH1GgEeivNi+7L1su6apFDQ725LZON4CWu
9SMAVNEkIXFD4uc2J8ikJDvlbs9pxqyfXfzRfltJMfYPypixB4Crje/TZ98I8TKEtVg3ZjDaThaQ
ygWuesMlES7/JPWONyu+IZ7wMuizAWaqW7PbGPrg91QfRpGmI5GWf5qN8phkCjaMtvyZC3WaDeFz
hph9r7DVb/ZCzz/7eLHdpPHxOxvRKQBZfzVcmFyaFFyMBC33QfA7HXUff+CluvB926gjpMVzF+89
jkELI6jE63x/jmNev51MmwzS9URKdx1Gxq2TRNdxuQCIg4hNUhAEsQ3IHarqsC4wyjZyBTOPQGUb
JPMBt/GNkGc1riX+/uPELF+ZBjG9PS3WLvH/XZ/B9ii7ilwzcpf5ekxJ1jmO8bh/DXx8z7qSLZi1
VLrh1cUZL4HHiGcGl9YxcKvINPrIaGJijLlgZjo2EnP8jMqn9bCGFK/HHLUyD7obE+Vk0YopIc2S
VYDRDVbtNPxygNyL3TVXe2tEntDT6vTPHFB/8c2BQZlxxJ9Osu2v1lYWz1E9qnDu5r85N/8mP7Rx
C9VnAXaxMIAUzruGnBL2mC89GbklDiysax+xI4Wb2G3G590cYBepFdL12tamdzZ1evSUgo3DKF4+
SWeG+81X9bxHGLujdcVGqaNjZigiL932U3L3tCT1TzjpI0tUv1yVtB3xt3owblVhT+7/G+Rg2WPd
i/RJVzqp9Xx2fApun+EY2Ur7ffxYqQvVmDBQ5f8DW7rSmd+IRgiJgPj1CR9h52Dy6KFpj9WZ0G0U
iLa7Kcz7Dz79Cyo1Fmz+r5ak8wNNZZNa8n5VDZwVu/QM7YXzvNsofYkzqyZ/XzIvXBEet/50BZZO
q4igz9VLnWPwuMr9DsG19wfgDOGAXCqqpSX0RFMWndvQBFwNhow9bqTKEZJAjf/GWK70WTnE2fPi
2ChDbPnfgGvBVgJtdflq0SYbxk9bXMfcM4JPaQMMOs3/qTJb4ql4k0qlKZRsPSa94Xc+U3/tYiDZ
esTKLraxGeW4jg65rtDHkO2kHQVG10PmIczVtHvmsLPjWW0w+ebBCvq+cWe+e9hzsE2+yxfMsy/Q
wTh0dznvc8RNKkIytF92KdKwTsZE5R6mf4kH2ZsFEqjIx+d8PeiFhksgbtS0DPSGs1jxbUdzTjF5
dESJ1yVUwPEV4PxpjWStpgpxzST4TUhYde0EaR8QuvRdlJXYkdtg/eD8sUTPGZZel1Kx8+A3RpNW
uqIhb9s5aD8rFKHRYr51tSHTiSDctfLUrLLVJQPRB1I5CVd/5az5lEyju0ipHv6H3RoXKjlwk62Z
SK2WaZXY4gyfF06Mz+A4mGCmxwSzTNnOdXGGBgURSg5/uzkrQ1aecOCaCPkBij+rLD0EoNDdiKVB
b0N/d1Q48t/WN9G6dXoC/XhfbxPgEsWvvHW5J+upOZdoZlru5f5+0tQdcBOMUdr7P0SkSKlR5UJC
WhBSwZ1t+zMrwDhHnAUeiBNCO7ExgAlckr+5ipJsewjvrNX4P9JgPGQmv9HhwAKo7TBsZ/er0Ju1
dAFxS7nWxNmG0Imw+P3lFFjirLuMQ1NDR5b6say71Ok54Aj5A3ogFYPiIcZJNct2Bq3SE7LH1Lp9
6BHyXL/WEQgttrZk+89dhNyQ97R5JXE1kF8vSVnYK8A7lqc4k3YKvnQ68mShwWWGNiUSKn5MGV8m
IB+zR01UQWBqy2ZFB9V/A6bA709WZ09xqIkDsbIMJqLZ26yjXUTfzbBgB0HKjwYzaiwoxe5bHBvG
05ClZDWInrL7x5Nb8/97H4laUcGTMaUSiZ7pPtz1WA9fbjIPw79NMRHiNu9gfQSBOcDBgf8YBVq+
wnvnaLYBem1AAbg9SQWrQa+TWg1Tw4YOJvY/ZPYmNg5eI6gp7It0K/5BPQgNbsgQaw6JqktmLuEl
svlWzv50cKw35RENI6FPsBgbU9bODvrqetkFoGjEi5C6jwkIjX5mcTfAXOzzO5pF9HKqv8GOLg2T
4n3JjnpkCc5IzirFFfsqP9ATZV059FjuuQ1tZF15cAsxUHtHWJiP5TxWnCrSa2psNaHw1ZHtts96
VHLWLGrv8IvS5wtP/u2nEyzZjkb2K4Tk/w22Ms0x8050EXbCv2V0E7W0yCL3mHr3rH+XHpAdqVCw
C2WiB7HvdeNGMt+96Z36xLvnw+FL26s4vReByHkl5YLtUcABcI1lLYtrJwks+FVgIb2pIUUAQStw
AzsWUR7bjkm36Yj3S2HhvJvTj8UuUamGZoe0e/aUVYKk3Uja+QcGO7SeZh0jP6FIb4FknSY1D0KS
n0pOik9btApJvP7B56iB0/o5hm+0EUl8k75YOQG4deH8Bf/M/p8FzWx+260jLiyOFEqmUTjfX+qp
SO6QfFRHeEQn6wIyihY3Td4GHfq6wW4omuDiziuJQ042w843FM7ATXOZZHaKJ905hBIAhKW26suO
OC/EHioDhje7OjgorWrwWMe3w7OSIo9yoqsFnczjX5KOpcb42dL9ujUgYfc4P1YiIY7tzpa37CIL
biGBBrACxa5dcdLIBVMSfRuiNfq1UWVzI6R2aQts0JjD2IzmfD7XUKgCSIlh5ZHsLjPX0HpKrnww
2JI+g5YWcNFZpdA4uZQFpyrbCHL+AYuXT8MF1tjcyFwgkHqGxRY5sGjEUDxTsdkUculWcA96C7Lm
UDSxHlgtZ0Zdv0RtQI26vr8UgggFJXwVQ5Otm/ccTdNVQ6PvR5cGCyqTTsMq9d/5JwQnkX7Fjpam
zsW6RCWp001b5a3k0iXMteMEFH882Z4OtvAJ9+Zq8/aSMzW+UWQ5DmXbLd5H5rEv20tSOhz3GcgY
cRmDTuCteimYuD9pLtTJpRXN7RFPD6WJUMelPsLqyBj+c49cPWOEYRNcCU8X5/WZk8fhZAIIxpT0
mDeogwcM+JMogxDEIPv/Kgrz2oFkyIBnq30pfDjqR5eZhmY2vW5mDlnDrZNV9vVuASEEo7VCUHx3
/tB/s8v3hUjVoV2p80s/cAqqNHsR6z9XcF4CRgJbqrFUYgZ6J5fmen7PuC87NBI3f3EkwCyxSw16
7/giXiYHk3xcMcAQBPDk6hB2vINyOBuIUYOJcqL2hfwqT7NocJwF1eOhXcFSqh9fhXkJow6j/28Q
yQkIuly0AWrjpaK8jTuwIZhJx77+MKHQTAjVKbPSfElLmZ+Yhi+hiAfX4t/Q1xh1ZTlY4Gjcs1J2
CbCsf2D9AugNfnt9HvdNOLeKMIRG63j/AwuRyeFSLXee/xUGjljf1trJlRdGqCFpGnzg0dSXAuIf
gts5H9cNNIWoSuTfl+jQEoR+QSmnVX28+9xC7n+JcXBTm9QifKzdBoCUYA3im1NA7nOT0DZDvAYd
4nZ+6/ZhIH4283YXUprVGIT4uiTe7HpbSi8v17dGkljZcHw031SUwDlEdcsb56unTxADOUsvfjEC
y8Yr89ky+uZsDEgoyZC47C88nVvtBm0Zk/uossGUSP1+d96+4lPn7tuEf7ejLY2y+Nn8neKFDOeH
Hh/O0gVIrJz/rdT7ylFSYMjPKWZKrn+mdip+kcmTv+JH1yfD0GCh+DLhdO+teWNoBjRHfnMIeQLR
EKKBpdJppvGSrPLz4+QndYOEiR/JAlLBQTgXmibCpJGZgPXKgkq7RQd2XfT592/OwrUkD7LmIIHc
jTQvvu/Ht2ouaeVDSMPlwBvlJPpU0fiIr512GfYc06qTDlWjQODw9JeffUN56S/EtLOI3rWhvOwv
/jCOUQrNmk3ur8ji/7BMyH4bkPhsScEg2CjekNn5YAFfVF4TzO4NzBw1ZVxTTHZ9TGcQHVEpqPlu
buNlhCDxQahIEaERufKvy/Y50aPkzpXbQXr0eewg6n2ShaHLCwJpfhaYVDjXO+WJ0gdgjg1SHnEa
ARxYmSsnT3G3cYDKAz6CUkVzcr5WUXSgQ1KYFgtI5LQubsxu7wTQ8e/94xl0zVG8HR8jHLnWnnRJ
9OGUDNZ1V1s5PZdmW4XGcNluv7+/IVrrpzGjahW+q/ETTlMvZlsbMGSjjtekp8JQzSD4sV9QP0uP
TCPD2aIwZRZMLk3L7hPDXm73vTeQfZrFwTJsSRwbenMO9vQ4/2tXOXldR4suxouDh7x0p2NNs3xS
2B0qobySPYvX8nSMJRPrci/47bm8PCXRnXV5t2iSooSVxepNFMOSqVm5OB/U3lwLtuELxTy4EmYV
1nkgoDkOo5/NjPUTYU283Fm5KjOunSzqbNdmjmQKW85LSxXI0Iq3ufCLHwchjMdgYBKZzgR8/ENQ
dRJqJerTbXVOSSGhSuCikZy5DauWx84iB3z4bN8I54YbIhcEIrp0o95EWm6txbspgWT+jDMpp6jr
WxJbKv7hZTngMnqtozOB+Vd4BudsxG87KK7hjUcNhIO33lgwwafprcw7szJsZUPX5dfKOG5+r0+p
sbOJin3GYxOvLPY9M7UHcDBJNjAfcnykSINzExxbvY2oN21TXYgZJZ9S6Ba7FjBuki8cxNm0OtI0
v7GGxEpxMFWJN6IDxtqVdELEjpo/0DFmsE2FXjP9xrwphNn3Fy3S7CVBFVM7kBcSYp+clumL8Jrq
lBOOiF8pWJMVfUyEIBv1m3vxsspZKpHncaEq9weIo4uGi0TgtLF1nz6DrVoaUPUhGYPnqIW/FLrr
jKpDfCPIcoLbhTksFouiihCLkAwqYMby6Y/Zo8aJ/5WWgWLNMhBNsnvDA37df+2+GGQTdNFfSwSS
wjTrw1RBVA0+JCH6qORu/hw3MW7sQ1edS6Fn/rpqGEBUEK185eTf2pW5wVGqwFNrUAhKVPGo8X5p
9OYRvGopnf3PkkEoPvVWO4tUein1R/xdNSrfSKHzi/A9LwYzOIGPUGaoD+YinngqsF2qSyChGzmi
hEXPFfEAXJzK9Ss7cN68dB48dJ77mKpPk84WbPJgBfVGcr/iNRAop3qIGMtRepT/GOYAwUk7D8eT
ER8swGpMIYzF3yIbwri67mDk16NRvTBNI2+0X1TFeoeQ+S1DLHYlIichFCix2WnYnFE4t8SemX23
GGXLT2J5lOWKiUgaWzui1OiXj3W9wWLPJn77ooMDE5jGreWlA6aMcXHz72O7NC+zqG87xg+ZS5RN
ecwec2/+6D/Ob5L0K9K4Y0x+KzzSKx6iNSZfOeR0GCM1mP53d19gmQlrj4LYt0ReZJ2PXl9w+1TH
GA2zL3Fye0wj6z+1Q4bQy6fpaww82o+cItfwik2tN2X0aDC193aoQ62NYJudpIdI45vFdkm80Ycn
ADLruADkGOCcEMUTlaa6xXZpN3/yW9BuCrJJaKM4OMoGASXzKv1ul1fqTkNLgzFKrOG0Ejz8V/kq
S9Sn61zQkVQq1QLVfRktohS602BMowFyQLixzypzLrRgSOWOAme1RgfpnFO+zA5mBtvGk6hxZgXP
ygBHFg6tf2BAfHrRK9gZSoFCWOKhos2j3xc3DsJeHdcBVyEfdUmXuroq5YZIlZe0/GGlBhjh4DEb
uYuAwaDBGugX2wdy/mmRtWFyd9i+YLQbSFpE+dWJcmytPs5Q/9TJGXk7IiQW8xkFszelHTE6iIda
sfZCTyfgOXKUFnv+OsYIe/J9IuMFVbewWTxKgNPLHtli0pw+46x2DL7wWBlCSdovHrzkUHzSYQWi
TS0CK27nCKohzfB2M1DwMSJnWSj/2EM+OVWl6s4nAj3Mot6hx9aYjv2g8Pm9hexwfXvTynIB8IAg
oV2vCxmp1xCu44GGr1Y3/JQ5l5j2QfCX2nw4h0GwkVLMO6peiHYtl+wXML0lqTn7vYOfUapQ/GK7
1zJNfJ8mo5s+YKux8FQmPQS/vl8aUPkck6/pIqgwGwK0A35WJA/3sFmvJiTphWynJZAkJjChh7IA
JPZbrhDzaf21Yo2lOh/AQsfabiaZaU8hScuSkJYyT+7QECgXTvnUeo9OWQSrDawDaIHM0kPNSPgc
V4fxpzl9LlcAX4cwuGmO7IeJjRtkP7e4s0SjNAuDipgRIJD0/TUTaupyKP+e6W1KR6xN7v+gunuK
e+vnwfVqsVZA6yV25jhSvhUJBX5/49pb6i9wLxBBkaPpxXS9Phuaci9F3qrLAxEjg6a1q/7edHZR
o/N0lkgrgFP7ZRfhjbj0Knt17tTDpXuP9pmiFlZAh7UMA+vzrDvRFHsY7eaOy4ZHMemwpG5T6F1D
Z05t8VOg84wGj1dAIiZmtzqKPQr3MXHISh8yTOR/D4HMQF4HILLjq9bZXjWq5Kgg5rITT5sIL4+V
omh2BX+Sl0R/6s61nrdIjNLko/PJWF4a/Jl5sEmD8we7kJRoPjGpm6EBDItkhBg7iieN6YNIL8bZ
aihbobNt4IiUH0LHDD+bBCvOBT5PJlmNkhhMe3x5IaDMsWcRoQh/XMIB7wPqCmpPx39wycOdM3PU
w1zNay/EuGB2OkeiIGi4xmJd0WjNvC0cCSyM9mE9bd35g6mjzq8K8RNDQUwhcnpDkv1JFAqWmssM
O5D4AWjP7XNGNAxz4a9W7qlgme8dZfFfiG76t0lYxAyM14GxdmX/byKMBLHuMr3/eVtoC5fjJxTM
9T3Bos16heX9xScXZ+MIEUHrImvPEMGsPsaq2l9dR9oiWGicMhcBMlsQ+/d8qFtFiIASRwtd36zi
dsEh4yJ4CvITqrUrdeCmr5Cg417KiKdlO7wtFV5Sgnk+PHvlMbIhbR9z8hnkrTEwRQNTnzgYYTiM
W5v6MnQIuP1hAaSpuXexEadJuggSsVt5xb6WQ2f9aKgieYnSydWeSuvqDH6NYM1zQattyhS4SHDb
M8i1EZ0LeNj6jQmlB4buUeC7qqzGsoChCfSL7jc3JfJ/tDivFmLCu2BnBZUvprd/WmjP1vV0gIB4
jghFmf3zNEsQHW+tS6O1yGsaqdiVdc4U8TDHJEVrA3oXMXBGKX/9vqC65CplBzMZfmYmO2aKjl0V
yD54v6TpFqTh2vr/SZdGBJAdJYJV59K4CAC+/nigqm5WPDIlAM9jC8OCk6D1i8AEwBJlkD9F5a8g
jxSai11a4pASBXPzkcCE2fsjairopWmdCQt+zPXIyBRXdgT8q+bOTqUcfCA88oDP/Dejw2N3cWIT
t9AyG1UT8JyhZvrMWxR9aCFzOUNDanro7DOe5WbCZYo+3V1cegKTrmSbUXWvEB2DIPMLZAyrKIb7
CPlbl/I3FPle8HvXQ+/jLKGsmRthe6O5KkgZNGHiB+ajpyZuGyn07JXhUUxR/5n5KPFOD+Y1xyTT
gsNGCMUu7MvHnY/f/3tPVfYysztBlnWbSRa81oFeXrN3y1PwH0dCeOFdJa+Uh1PjeTQF6D6vEt+V
bVd4iaZ1WqsULqLdP8Oz4vXO2cEk0VWyHTUUxPHdGJms7cldLuhz1rnx3JSlFprCOnUM7NQl8UO6
G1bVr6ySiznW5NEYFZzT6MoujQbzD8ix7e5qXsCNoYyVqaE88fWaaYb4fK9PE8CkEynCzkQX/cSx
kOT+0DnB8UZ7YyYD7AwOVTGullfsyNs5X2NxT+t5+MqVnYuAfq/vqujF1k0/jw+JCQ0gJnrPIr9H
Joet2c8I15wh/DYG3SxmZZFj+yeXZ3StDm5/6c+aDW2CfIiv8/Ho9pneuLc3uM8/XXCKLPTJoDTM
dMwp5dI+LJN4QbsmH5Rnk6DidowUoEvghJ4gxrk2PtQza0ypcCejQMip8+A25d/M8CtGNYmVgN0M
1YJdu280OMspX2gzwF04oJRxrjKZDYFIJB39VcgFp0UxUhgY/CFG8TXUAWAJgaeE7TAFvGX42Xiw
20x61OoDh8l1kzUOuKmGKW7sLunY8X+VAJlKh3OfHrFPHpyBJR75kxKy7sciVZ3a8h/U9mTiyP8b
arjk/w9j41UaieMUhmPexMOSSFkGZd56Cn9psM5xG3RahTUlVZVaF44jGL+Xb2rpbxBANh26N3hy
arhPdQ0qZ8LAFg/5cp5IZx5rpUQ8fIazMK3RNsa0YHgEMMq9SPWbGdLtX5dBHK7FzYRy1bD0+C6d
s90b5N2Ae8m8jeeDWFXVy7BQTvWCVROqqKx2UXNJdO21X17UiltyTywxVVHlIIhuTi5ynD/R315f
pWKh4jhhlx52iCpthBmyIhx7GXDebbsWC5hdRqWw9uNhCDy8f4usgpepNtP+tsooy4hcSNjmL8Wf
71hf8IymGWrtCeXwfwsj2UUQ4HWo1q+rFnw0n3VqGWImUvBN1MMoFW5xGZ+xziQ/OAB+2P07Ns5C
uKDpeS9wSgnPsC18nrMjDa9Sol7BlTKsJLnJ8hW89d63KW4bQcTkyeqFuEOjjmZm8sg3qahjGQqG
hpCvKj+c+SbjF9ANw3L/HnXTdF2j9WXoj7ErgGIPd2VP3ZQs6YwEEaEXK15HHJe7a4xsXAiLW+7J
zo8lVwi7EzYpwz0LhFgeUeiMYyiP1bqMt7jeH1WJjuiSTcQ3D0ulKs71Vd0tNeQ1T4ccN3QRIOwf
LO1NFjWySKRrVlaPODeeyCZpRrWmyOjeV8a9fPINw96IyClWqMzVnYwSqlJ+zOSEtTmDHoFit2Fo
mtwk4OQkU1cVeyCAYQcR/NT1PTRk8bGbVxVxLUIDA+uf9BoawzrGoMtta9TsOWMSHA192AQtW32D
ZbBuMGaFSqL6Gmwo6emSXykmD52mOBHn2FEyA2yBq9/qxb7ltwFwSnlja6UfdfNfsaFPWUusXAFp
tvqd7UQ9SlE/URD8UGjRHrQt1DDTt/QJ/5xzcB03raH0gCZ7fw/M2KZLjM4uBrvzlsYRE1jQX+8l
arnwnUt4kDXKvs+FNJcrL4ml+3hIF6YUx82OspVcXfcxSfeOje8iPv+efeXUWWkPkW19Va4lp7Wz
v4QTGSbVdUfeSFuknBb3XascFV9sRD7wLCl5oCiPfzBpqgf/2/DSTPHV9AimsHrjGx329chRQMcZ
Kgp22/SNBfterOaoeww7pKtnWpmtq8poz9TEJ2Fx95E42LlXHB37Y8AFQ1XbMboSkYEQbJ9XFF72
9fQqHEg6GhFoQp9uEiwxMQDCWJUhLbOC0kihXRXEKR7FTRa6XtEidXT+hQ/PAJA+XESZ2jrakDZs
piEQg6ZqTwbAHDV7pa9JFAULAb0U+uBa00OBvI/pEJMqagq5llYZYbFZNbo0Zs8HF423NbDx5j4/
Uvth+TNp5g2/KApsmSgQ97XEiJSI+KJPth548gwg/AQJ6tsk5YFUMHI4rmvitf/HzEWEQLgnWqpe
8wCtpx9E4HiBGRtkyLWPaJvLFwEr/Rc/mH3LjavezmhJ5qTN4VNAWX41YFdVVa/ao2HS5SqjNAMh
fnOqFYmsulOqTzoRpfSqZA7u2ZnATOU1ix1xlKSsmdxow8K5J/tOp+f5VAlYDuvUcy90xeLRVbTO
uzV0VhxHcdWHClN0sG/HV6h+ozTP6xKetxK2elZPofDlxY1lfeiB6LdiNMkT9GAsSoZSUCSGVtv8
b77z2L1at50XdrNJ0OfTVSw5gaGqZm0dLi5bZ5ukcV3uPDfacqRmUpqCcLxZEG0fHT8cPr4082x0
GAJcItzP+QUUlVpIXxlJJbvycvvjlnr1OTmNjTg79gMGtUQD8WH8AcuGXPTcX6YvsOx1aSsx36H7
yW3PcknbamQiowjU6bUILXyHvcBBas6BixrYFliTn8r2abZxtsCStYNR+Aa5oGwI/GUMYdHUHuzy
HHDTT7kwHSESuljTf+62uUHuqSWvljWKlJb6cnP093PUM7QbLYTXVWpTSRyrUox/eatJRk/tBJ4f
+LlRlR3YXkubhj/26Jc/4TPtUZ+KezLExi4PQCve2lFdQPfrA9oZ1JYSFJwprt+U9AkUvvUlj2Uh
R72pXp58gS2WSU7vBFqQCz9zwjEnKoqqrdrMoMphQaXyvaRni8a1MOXE0RaeDYfZ9HCWpTfWtO8J
eXpoMW9YbWr1EbHdrjWp4g3EQ31foOQnHyq3KWB1KxdHT6JxksOg9fAaXUFjgl6H+qxCk9HeQXYr
RqSkrC3Tsd/2nDhjAJ78b7CsWB2vtK2F+dvLxpJ4ebNVEoUG7mfs2jtLnW0lt6B78iNOvMC+djgj
gAH78NmAUE2InV2k0AjR6+Y0qigx8ffLp0vGi3GAbs0N1BcxwEnZ9h8qtTWMdccrUy8t2rGuAFgU
rLnApGCinW4c7zSiVQdjUa96PpbZp57kgDuWCUhQtCvB+w4eJ8nwdZ7D25bPChugeqVHPKC4MfPY
J77WSiJaf1+QzlxQFyPsnLsxjzc2H5Y3Cx2fqKmPJQ/fJbEHJFml5TsO1Eo4bhl4P0ZktAJtP0k+
ZRs++mcZkmx1eKNxVlkzZxj9U84ItS0kKVvszAGX8ItAZhgdZsFymQ9TusNb8vmZHEQt3UZbp3U4
e5oLn1wEPEYfGpao3eerKB2KbfrJwTTD2xwncJv7KFD+8pDIcFLicLIL/np6xnOij6q23bUX5GBY
D1++Vi6ZiBP3r7TqWOv/ifIUWEGuI5w43BotJE6Bd68AqpcWluhElKzL3z60SFY7RINCfZrK0v7G
P92lwIjS4/UnSnj7Kdv5Wy4trRurQxYV7v8LuVihe+ezas0RbVl42ZwzZZhwGq4mOxVpo4MysxSg
bOAWkC5UoatGn/Ussj3kQKR7VW5WXS8vYa18kNm0gcziT7elwzly5A207EeSSHrbkKen4GPdTwfS
PUQaWNjeGOxZWV9Iq82hSY+wgFWbW9Qmf28lCCZkscBMjdxmmUXOhFYlE7VTSRVvgztQsy/NIGDw
UK0K/bXLb4fHyRuz17VajpLgh/1iTBD9F43QLThT2ZEuPgak5/bcwEJjNl+yAko3QvYGZ7mt0p4K
qcxbQVK/yURCDh0ynkeV+ldS1X/Hgk1dkhJkqLLMBwPxEvsQGCBPkoSlKglK05+h89grmaFRjigz
Lmdde2x1fufG8CnrQYXzPL0dySA8U7450f5VECrsjGFFywRnZN5nUpHNLwJOB0zLHkT6Q9VLZzyR
oDJUwwmL60kRNV89Flukyka4k0v+LuuutYzRClFIReFH+iiEdryVdIbHSz6BzgGrQbgVZsmZhs4J
6uabOy3RP0z6JOXSh0AJoqlVT80DxOLBgb4kGjKvsnGxy1RbnG6mg4NJhP9UWdNDbPVaqMSrHS6R
ER9i0asI0f2sO02TJNZZA6n61rSv3k1Ml2ue0lHiUsYLYOMELGw0juJU42G/68eIzFYPFgEItpL/
Hi3Ortgy9c7A3vw5l0TA15Q3QrqAZdW78BNDcLjQKxAI4edvVNr7hxr8FWTShH7sD2GvbI1wVr+j
FdqSnSpHL31aeh0WjzzaiGrMgj6o9j/MzBEIByDQLlRhPQdj3gcvjejbTlna6fKDC+5fHecArbn6
SjzDuxvMocT75PaUD7fBX+PKt0299MwG6/VG3pIeVtl2ZkL5FDZn5BA/4WUu92OpNxsMCZKQHvnS
EARG78UrEl4XrO91lLBRwm9bF14jZxAB2GX9jng6ExT0ZqVPjyfNVWp18G8vZBwGFPAvlbi0Yiyy
ZVh9xWk5VJhHICMIhEkd1hl2foS2fEJg3rK5YNjkJ50N6stgBx7UQYo26CLCqbfL200rYHm9uXp2
5UNA4b8iSccKuLDhVo7Jm2rYIhwnFgv/LnaAtwzhytwXqPNTFJPd7hn00i1JZ8/MABTsO0LTu6ea
cU/YHI/z5NMojF8a05nWpsVBpQfpSMQ5wwBpP2UPKIuBRlYy+LgM4vAH7KiaYcEhYMw54dVTpVCm
gZbg8PduZ0yfX8NMRMGsMQRYY9Is2HXjb4jMV3DNVl64k8flD/sJmE5BsmnpIYvMdVAUdGn5ECKx
RiZWvFQ9YZ8wvmuveiePLD50rJ/CjdzOdUX04StN1GjqXiRDuJL2txR5km5B3F+3aGjsFzgUTe9p
526rmziNMGK0JVpah1qvMz+9ZPSDqqiW0FcYBz2MhtocACf0Z+D8xf5Uu/9D+o7TvR3TBV9wgYaT
MfbNRSGt1yTJMyvBbUS75HCjuWZYKQYosmU+vS+BiE7rZS1worg3DR6UdCOyixH6dDdejcE61aSt
CH8wauu5NtUvYdQXWZDRRRbC6WI4DmAa3rwPWJ/dF3jV79XRrqj1JQApKiINiyIhxcwxudVRLZVo
YDfDXConwrrj9z9TpD+/ozNkHw5GDfd4NuUPuK/gcL259FLDUDx3e1YMSOuBY/EeOcd0ylTKIqGE
K9biTaCR7vbHUjeYv+xnSPBb+33Vm7vDijtj++hnEMyPbZpFy6xpYl/oI+Ct3t0j08a8H4cSLik7
IrsFvlGJ8IQbxQG8fwrZ4C/PGs4sWRSomRTSh3z0OidY2CIoaMXtuorPvBs/v6DYGSUftwu2iMR1
vVsj1Lup5xq+8j6REyPsJ8667X0CqUEodMAMEtvUsD0qPJJhJdn0/iQcDxhG/SlifXIz+YyKkYsf
IS2Ova+vNBdf/q0E2Xn83AAuW6My9vswFBvmG6BUcwF4mEX2C8I8LyDVMlm4RZtseYnjNswovMsy
BWCP+JlIuv014AE7qI8jr1RfYcbX942/1ir61xRCMMn3JjbkJA9WSN6T9YCO3R3K4xXvZOAble25
64Mj3zKP8vU5BqVLoakHlkeNsl1Rw/zcYEwtI+oQUU8Gl8uBQ3696Vw1mpEKwKShu/7iuzAhkUD+
3gl5QWBGvs34X2UEh3QhN1EUQ7Q0TrKoASJOh4m8Fu8wNmcicwkg8FDRldZ7w00IYH2TYaowhHxb
1S9XAyjPGZKHlKPIfELGBIJzxtlPnUjDA5wLTnk2AqttwlsKtNviU3pjEt21OC7us/l09KoxPflT
r/OEk7JPEauzL4UWs8Fs2mgcM4xKJ8ApwGm+2rHStSdveRamwjAX2higxT+TLeX0xschBiSIx/qn
YafCdU0TDBQS995z6Hy2hSgeR83MMgdGV9UvpM75PqImE1yaBEgJNu7RB5OpzUMleGT/h52/IJ2O
zYWafHRZ7XJ22SIWOaIcx8OlaCYxrcGHb/W+78bAWCc8/0u4jiZ/B4rxQUgbH1acjrI7Pgfhl7ZR
Y6F+WoJcPzza8eVabmvY5+ODrpeFNSLTCurpjkpYGffO+1DHYbzDSFTYnel9rXFVS/rggubsXAZI
dTrvP59BEJUodcHyWckFiixOcH8lFqvECDuFeeG6sT0+n1VRklJisps5zBf0sYP5yOlRx56wSCn5
HthPOJ9hUgC80sDZQ7sQnuEa9mTv43VZJfyO4Ovt2IXCTuALD6NMUDH2gWBOLI4naHryQeBUG0lS
W5quC/nupOoF5RA2iz/U4w0TGTF1TN5lHmgTQXWIAIQzBtogMebH77aZQLXajdOtFMwdAK2+8trh
/XLEZl5oXjW4Z5u76O4wq5znovoGaSEDoHsIE0t74OUFJi1GVYWDPvH5lUBoQMni/UXezF0vH1+r
TeNQcay8WWvfkhyti+5pA7vOI6iRmcXPDnWagL5sAnb7pQcI5i+3EKhp6fLlo7Fbq50GL4Q1UR6I
B47jLM034gigQ6h91A6RstOjX5/JFdRJHHHuay338m++F3jedgy9/gPHpgMh6K3dpBOdcHZo3aWk
X1Zlnc9L9mTvoYII0ITF6lRzXdJ8ec1sXqnSOH5DN/w2JJQi0dHo8mS/zB3g1/NvvfvgP9/t8r84
Srss+U0b8635h/sC8nqvTA4y4euUXzeC9jc98ZoEVqqbCcaAz4T6n1rSk+J2uzU2FFuVQelw255O
Elz+waNItrrUZiXXkj0TLCtSgMOVamJZQN7ONZVjg3L53QVogXs/bytexNrI/NdWpAgS2oAR8Egq
uWcYrJwDl6YX0YHzk06KmQApIS/In5idfNaeRLRAX/DM6+DVA1EEugL6aslnGWb5OWj5ysukTiB3
nY/kXE1qZWR/N3DTT8g+/KE9uZ9/MB74x/w7WuSCBtgkKXRGyoL5BpGq0dvEVyufnesPeUGdxQl2
uC14IiLdGagmSsWEcGWrbxS0JZ87pwrUIQAj+9BeZnkvB5LcRi0Ab0rt3ZnMdOuXQe++q8J+4Hf5
pCQJe2/rhp3F386FxLFySicnfFvWB9F6iaHCaX1kOv+rquUXj2lwnX4cz7FMGtqS2gQIkvqyC3BC
y5zngcDqI0hzIglwkQztv+1MGeTxhlTy+O+uAy2icLiNLFxq+XM4LNgAOaRHsQcerrRN0v5SUROH
6/du1r8++Gx3kEluhxuSkr2pxtpBtgVOAQkhyRdvF1y9xrOi+OueBdGiZCN/rywi+w1xqiWMqf2u
waBWvjjspbVu7uFaEEU+Ji6uUKi4U1tsX7kog6MWOGNOtkZFcKvjNpwdeJIvmBBXAjB3hT4W3pMr
IjXHvZgzJ78ONB4jKF51LAUl7+pmUwHp4rBAp2X+bNdfEXujJ0HqmvhihiFryotp8JazagQClwJs
bTH0Qgr12ZM6yWZp6OAkapiPUuvZE/B8WMEByFJIbx+O55JZjsIVx3uBPmtkhRWkeKXWgmuYAovK
0y++HM0Wj+1yErn4L3pMTquI5WtY7jHJduCP6M9GZS4o2jbumBP8GJv17Eukp+tyRdVsqpclBJRd
6GKjC1q0JAo4y8Gyby28Tn/Z917ziMjy44gXl6hku48ccqAD2/jWChKkyJ5I6c2V1cn8RXRPICK/
8BiJ71J1tAB6WAO+333etSQIpVeaeSQSiVFG0E13YDiTfkHrvStSvBuNPrfSs5Vv9gIu/qPeUrNy
KGgOim+CZpOhAAGbB6F/xnpVFgCbUBmZdHU1CQ4j4NxsyRIcPk12JfPqIRoioNFdyd9we4NXb74b
mE6HR0yrdbAkTBMu9CCFn/8OkG/8wVGXKaFcKzatQJMvNp7Nxy/1EorVWXwLalGtVQsgX3l/6q5p
CDr7W21AzhEJ1KB5qlxeHxpnR/lae3zrhclcBF9ct6H09yvjwtTB8trYYWhl3JgfNZJR+qIRSY0q
k9XKCBPgtLzyL2PN5B9y5obpf2DVQ2O9fO/k/WXMaticAEnrbHBTwRymCzf90EWIlUn3NNjIYePB
3gJj4HtoMk05270ck5X3x/m3u51wCckSxaLc1dVyENZiLZhe0k7QyJ/eo23mgEGtEeK42g+JgT/2
9sQ0wMKgdrgYQFMHXzKOqF1yxUOYKQNFsfzZDIQ8sFoMhdheOmFMAkVP28XIQPobI0slSjCeaoZn
IzHpLw4ZFX2wjo2S2x0fLWQuTW76Do6YAnMjHu9RYa7rZ8ytLZYoVzMtWHYu6iddIhDYhWhRNhiV
2AFMSN0ONO+BV42+COVyRDh4qRC/i8uDj7RCZHcLlfWGMujqC+WLQzoCs7Gf27sQUt6uzqlhtMam
3xDoMYBH9MYqYo2RfyNiSDyJFnlTwE6nwILsIBaLV37ZDMOolCED/sf0TGHmbTt+QRng4bL023YC
bSJBVVqRrLtmhBeTJXoCxDiEsH2i7ULL0YuGAuscHDGjaz0qUB6yb3PDQxrpsXcl82I1mn7Fd0wu
4vyB0HYD25erIhbZsemNiW5MIWxiBtoNR3G7mbhTSda4miL7J4YkBG8oCBc2shHSjWmMxgWTxsne
Ly/kEaxcZc5ZvcI0bHis37ZlFqYWmKgOnA/jx3dbhUm6wBCCKuryVTs83ugLa5vzPs2ESOcsNyvE
o0OHY7ZGsn+D5gI8beLq/JPNj41k9ky0A54BP1bs3NK4UIDGB3LGrjQTy6E+geYQ5ix4f7fh95k1
tn1cS147bkcdy+ZdVQx550AOi5kolFDQN/jFmA2vH2Ya587M9kZejJiC92Gi3HQQqXYCb3RwYpMU
abgUEtuAdYakPVOskI9VljdxI3g4SPAX0fzk21oLDldERBaUv0rS5ZR7XijdynjpvVkruDCBOfGe
iIRiQl+g5sai/mhZ4YvKCgF65cLGyCknKD/jhSxP4jC3bMc0eNq8gbr0AHG6NyWGd1EK+RXpKNDb
epwgGmvjv5QpERUjNgLBXBNyWVES9RXfhbYlTsyiuQjWG4eNZrInPSE06ggktpjDJr9t6h3JGZJD
fnUfCjzDpcOjuC/KYv52mt8ZdKkQzbgRpCVjHxMxCRMz6Zl6+h1LYCIaoMmk+S8u32JV/fhnKAiz
Kil8fW7vi9caBI06/jC1iiAXzBvxiuv2iprr7+9BBLUmm0VI2YbFZ9eQmb9O6eEhqGYT0i6eZmki
/agVg2v3tw83HzsuhBp3E9s7dSvqxxrWvEMo8Zg1Erti1KPlHeveLerCdHq/yguJLu5p7A2G+RCH
0Yfme7YtpcZr6W/Ng2DqOk4Tk4h6BYWOwpiqy7hT9sel9SRSKNIOGgs+A6C1uL5KKQnipH7aaHeA
4vbQ6VO48NInpHz9/jtaa6RsJuVH3aU1lGh6G2fRZkDWB99r8Cd5Yy7W1UDC+ermtW8vRXzAbhC9
x2R3/6fkthmS2zSo2SVdCYX7LDO46z2gZZ0P/vrFqqmB9f+VjwlDE0pAzFq9MB8JCtNlPgqBx3Dx
OzmBZhmf5Ae21Ox05/B05zkTf839/BNsOmlCXzq0wS2HlGibkald84j+iB5jrWwlPts/mdR1VtOp
1Ot5cJl9v4EbdnINxw0usvri+UAnf2fTPKXL09j0YryMm1seopWdwzwO8T0t9YIcAVlVzB/A2H+a
Rjk7GObEF5Ore1EOqKlNYWxs9WdLE0ROanPXixvK4eB/0RKp1T64zpvnMgVK3F7Q9JM33WDDuIHz
yb5VSklT4hgq2kugCSV1boaOLAQmlVdm9ndJaIymuN2vJCNvD897OdqRJjzfEIGbF2kz20p0ZuG8
CYOcQ3SH0ODySbpB2dGA2Ppqy8YM8S2GMyM9AtKT4D24C+Nv7gf8ihbFI3elWn2kw8laCi4dlnuM
UuZ0NcXr1sUzfYPtCfrmqOrH939Jw2n35vBv7NWh7dMASfJRhUtomcmcfCkv07oi58HpNiGPVt6U
h86dLu39TULSvRJVkF5YT4JH2Zxshf0FA3ErDt3D6+OSiInQhasgnd4kBixfwa3X1IE+Ku0S7xng
qjtE9Prb86ZfPh9USIPfU6Fq+KJk7s+m1lh48E1IFRGpstTRxvuUGo0P3Suhip8lLRbObSGeGm0a
ydYgh1RbdV0B+lyKiPr4exut4CqVCcMcWl2+NmGivGDUbITEAsqJZpy4tqtL1Y/MRsWMSrN90NU9
LtLXacDL68wU79sB0ZZYAPL0j57gXnykqHvF+uL6GP75fkeVA2pDxWKgXFhYB7FqcSc7elohywWT
8s8w/EAVCfbUpBf2s0jLCumNxvyBy4unhEgLhSxsNxVJnWlHqvI2B2+NyoBF+gtkVeq5omT1nlmL
0F2n6hUGOzmmscdVX15LZqhkHHPyyc70gMVmJC2K7oxRkRzyR0BBhbLmkfMCdU86WzJ6WJNvHlG0
ZTmP0K3QpL072u9lztyhYLK1kqQWbdVvjCKxH56KlXX7gOvI5vuIlwpHbt6XVYHX2nmbAx09v9ny
PDQpCwdDFfwunDldJwgS8S+gxhiOIA2lpetCDNFUUUhqWbnm1HrkNWQtmMGsRUJGfaPalLI3fchG
rxwTll24TUyokyxRek9RPaKUxpp8VFwmmFNMRgznYaksifpzH1Ogn1zhjgCX0JP2YiziOSfDQ2S5
ockILrcnv8NdIr9y1SHVYeTcIIbolgJKBMKH34a5AuOZa2h5gnDk/TG4fdsox6as0VoUIo8h82Da
VeJb38+OVDHrqmvoqSGGGMi6ifvzy1OfAoixy3lDpLkxpCKXQSLVjfFaBEpMwsaSkweGOLtU+b2t
YIK4oFgwD0luLr2dX/8lYlkBiC89CH6Ye7/gb1ESYVFL378nnr4rcXit30Tqfc56OtY45jDBcniE
/cc4J9zrdphNjm5UhKZnT+MoInoANv/H316+wxj2wSLbHV4Hcqqr/1mwdb1K8akZbJG8cJOE1Mh7
qvU6tI3R1btD9u0/2Mr5OaGGQa9QhWO7z/USQUVD9jB6OJqojqNApJAq7ZrzZMsSnu60jCxEc9Dv
aj4Rxqoe3WO2KLGolAPky8FD6v0lCLxtOyzZzG0Mfar/WrV1tgp4DxQ0UnVivZya9yv0wgKiyW04
PT5SJoh2ZzLWBNVaPZIjD2fGkDoqPQ8qt4r1br48V+qwY/7NiOVZ6tWeRdRtb/DnzDBiIbNRd3dI
7wt16QGi53Mp6NPBD8b6/RY+hG7z1a2BhJvh90h3QNZh54tgtP/7S9V2JNwdWne/DFJj/YneIQoN
Ug/dkOVALo2NyrG1Qhr+zL/fKydv3VClgZDJvHHs6kdASQdfykdsB2jg28ZO+MKElRYAOdvKVxzb
fl5gZjg3OmC+mx4DkrsDJ4Tt/hRMsnsK9ZuKouVSvbFsGmcYiaPttGPj7Tzx7kFLvVv0UE/suAC8
gdFS7detJUJAlzSeFTMT4Q/wf+IZ+WbIdpQ8GNnyra5ZZyyHOvGtQyEAD2kafQKWmPjVSxxIDTkr
X90u8ruqWK7F6f/zxFfDzu2PnhC85usDsHuD4kvPYHXuQ90XaJXdiPM0mMKbNRv8xQpjB8vIM38Z
gf0CSWZuBO03emYzTBPz2J0o9zZC8mhyNYbOB/qugnHm2GWeizFxV+CpneeRQ5Bfm2FIuOCd3muf
hWFN7WHyCOWcwleqNFRqRm5aV6I+g0FOBpkVwlx4yKo3IU33XQf+f3s1/RUXIiqXnV7FcqVpIC0A
/TU2eZMWPpfoBSsCGs4cPKn0jFY3lNg5l2L4gAYAHNUwJQCGJgngNYVGu+Y4ZFBgZYFiiCLfSi37
F+aFXf99Iy2n/SzgRacHiABPul67bUfTUWEW5otqga8ibUNaFgLJd1dNF13rqrjtmx7NYZEr6Aqr
9uUwl4lL5JiaO+e+eNHStKuph0nLKsiIo0ATyOx9m7QlSNoRaKy0lfNBCt1wsmjhvvEti5iGhpcL
yVWG5HTpNGt4KEjRXhs/11O2gJB6EUR6PEEgrY5hJCwvvxV5trbpd0LQcS6RvPCDZXJW2oc7ob0h
ue8IkTvcP9YvhwcaZfqZp08wGnPKcFFiBCZUymY8+a4uvmL0DJ41OG+YjRVcNLCb15txVv8Z1axF
fZ6TNgjyZqQ/UO6RDKNC+iZNB9tSpoDpBvu3fgI3x4ghHfulNrmfarjLVSSg5BmP4ZKSxYkG3KX2
AiC94GkX3RxQcWi/43sCaLjURm7p+cY82mbF8xb6dGuFWgfIuJqPH3o3Hgh0LSDm807UinWTOl9a
+OaD9lfU7XTMougvMgVDDuzAZtXey52IbDrIomQWEH9KCza6UCFfrboEkRH5KXuLeux2r0OqA517
30fTLqnOghD98QdtCpxqJfp5g5Petp4qoeRYBTRFLzLDqWanFpHmYvv1LD5xnvJQyvXLyoTyPvzY
DVQztMI/j0s0QIAmB+Oe9PeMNfTMXm/TuTUbRkZiHGr5n2v4gtlKJf3sjawXiJYeuBzgVh0JuO6i
EA9eBnoEXnH6vr9PvNil5ORnxsicGlrTA8U0aoZdo4BYoy+ovxyaiEZfYLW/QqY8KtNCR5BuBQ1X
gfWopgnlUPUouwqR0Mrwc0BRBwaI/IWmrt8uB63BX7rzmb6pQCnxUV3CAfpimgghb778Q4p0F88+
+oaFbQbrllW/lDXHEVWNiFpaDHcBXBFZF1IczeI9CkLKuanyUyEOpGDgAOdIw3wbn9jdlg9oO2HW
YZf7Stxh2Bi0ryKa91j98MIoGoLUg7eVFYDjxRzgCVWMrh6k9sireqd9gBP55y95FCmrUladooES
yuiCKbrmc/bcs1P61dVJE361+gItSDWu2MyXHGPJqImtwYJlo2tNa8MR1Q7IhcWrW1BuPcZfTtzv
FC96ecAR24SvKi9q498tWrsLEptBbrkJnDPoK7NaSpm3LU67Z295JN4KrDp1mE75cAkjP6mTJY/N
F5b5dxnYM3ndD+N1hZoWHZrrJxWaiWLRo/ccl+T87ZU5roU+K/u5/MpCUza0nN29AJYnQVcrDQei
/H+VoPY3gm2eAX6wqA0Udihf/Rssnz5bcDoGMtFPODqlZ/rAj6WCvtHWGPixKOMnOlWhIgYqnl5I
xjkEus5l2H+UpbN8R4Hs4d3WhUBWLx4IBUoTPBYMo8nb2HlRS2bngV1vKjnJcBd3cdK9f9ZQUMDb
9WE6f0nez51NycOJuu8SJBZ2FNfSJks+ltI0z+bV+KFWAEwQB6JvYi5woaS6vaKG5Lz/wEPsJ3r+
8rA+LNmNTYGboWk3vQOLQjR1OSWme8IQIeHdhVXd3qzPbIjgDmbeMRXwQmmsDoPZGU8EMQLzDCL4
FbSXPwMARKeC61msVxqF+h1ETSQ0Wqf+3M9CnszK6psdQ/Pfn8n/G0Xlu8+QNxB2THhvnMpBZXPJ
mLO7sRZ53Q2dBYVK1/BNnsZsfVhLMLdqbI2FVUDG+0pT/LVWXDnHVyoQJFWjDHe6nIgsBgv98tgl
kgqeKzsE0zDcxC8PjATAyQ6W4ZqU4K0mgxRU7E2J/xzvCq/tT0LVO0b9MKO5bEWWXkCM4WurCcuO
ACVqXNLE1LpglFDK9+FqxBYXko8XYbKwE4Q+BrKNAAwzdS7H+jHqTRhQ1l2faFTe4EMytMPN1irK
IXJA+02r0ItIxEMWdEZlUavbFmeVr3+dHh7petJWZlQHpyD2Fy+u1fuItvJkuT+KguAhQMWzNsav
211z4ygh5sIF/Ypi4Ah288hq6jRMiTpFZiAP3N9638r6IACN1PApWzfDVlIwzwf9HXsH2ih1DyJw
i0t25BbpCFtOqsPy/8fwmFMpstd88vMRDW+Ka70JaQTPsjTvvt+5UqLIQ6xgJbE9sfahElvAch0S
4dN+5Xe9Nfox3/Zp8U8RcgmpYycJjkERazZJ7tV8I4AhYNrtJUmzW6OmsXfcVH7loSYHujZTvooK
372J1WWg5JvYRcpcHitrXoLwPTvp3bgLPSlzlkh5bw4ya9QrJ8+AliELVbz7pxNisScDR/ScJBtX
HHw3RXwVw4ueIAi3fzv1iSo+RtXKQcNpfyNQhbzaoo5fHB8voaP9YkydNodan4XdOWST8SjZFpNF
zt8wAaErXkDirIAAEFo9rAUpTfmh+or6s1+sXr5LIsv+vVQh3EDUWYcFFWEnf3oVaTe7a2egR0o4
gH1jGm+VZ7fv+G7yU4aL0m28I7D2OwDVUNUrDVn2kjQV7pWNFU/oz5S4LvQ90xpTpnETGIMOrhIE
fmjto8gGCu54M7VSG7C+jpe2/vfVB5r2HwYjmBxQbaBkLZD1/uOCBmtV1vz0i6yAF2xTVb1BQTCf
ZJd4k6/fWlKKyYARgIhemm1wy/qCeDtE79mf/RJrzhRWyYwx/JptN1JQ1cSxAyDdWSYka/FME18t
Ol5a3u7eUMnOT9Mdzjc57Tarcg019d4Q3h0WQltlfOaU6ZAhq1en3Icn4IM6UHWyLN/afrVIGvnB
vyU9hP3xzM4SjLfy0H1ijmTtoHxbUHDZttbLPSyR0DokLQ5MrIWjSjcpTSH7D/l76iaxmpe+6gkA
pyIlrQ4+oorwTB8/U7bkpBFXbtflNptwwevTR09MFlvk+YT/lwS37Lw/I0dPR5Dp4M15cAqUf4mL
mdQeqjaGK6nUwBV7sgxq/TnWOEfDp3zQeoOOmWbeXQ09wlWIVGLN20SVWNXXD2CIzZzghg8Stccb
H89qK9TS+7kmPYNbeLINpKt65693R3eeM0ws2zq7dRsHqxxSz4oouno4XrZnY3whEQqSze+nqMZR
rhbJRWl5IY7lS7g+WspywKAUX20XC3mpSV6YM/L2TW2DDjqJ/zJyYjQSIneN3KR9nGKO9pQOcKXV
ZFzbbTEBDt9id3hQ6esd9IKIL2JdibMyDiIVm3C9oQoXIgGsbBgYuMKe/S19h+F7rE8Fom2Vf7t6
DsPuWscoHvpgEcFUk7tA0HTDfMUAVCgnxGjsBLjnWp7sk+H55eF5e/NFyJmVHMzZDHKXe6DuebTD
SDm2yIJp/LkKfmcCunEFcGrOxOnsR2Cc+AQkfXRRT5KRlaVn5cUiROuq/8uVsDx5qQJYMDGTcCqG
7TWyZ8akj9gXQ6XPaELe9ll2ox81HHlQ02srNhlleWJLBAJC7HHgNaZLrAJaIchRIQbnyTHmGU5Y
xRTKZHDdpzjzEMkCi20fcBywX3ChZiBil8bKAgqNfCotLFPVg1pAqFGlG9TP6Ci7iArdcwAEPi+z
keysrsdH/VYR7exPuCXxtlrE25zcuSo1s6JBrc5QwRjXVCLn342ggs/ABl5DZZaGeaeCiH+ScaFq
+4A1gB8UTJcCMQGqirkCVRxk+M/N/Qr6jqIOcJtFz0yfPHfdn/GX19DDIqProBE13lipWmqceY7I
T5NqtQo3UEzXQtKjhrAFOK6zYcOAGnhNjIM1J8Ow7UJndvodyHtyaJCUoQd1yi6Mrp9kwAe/J8+2
02jOVuaxxlZagdHHtjmMZiJmMYwFGJ61aTJ3UbDMLoOxgQGz46gqvQl24EJw2XSuPhzbvZ/Jgu73
ElP+YnldzJBVVGXLshe7AhaCiQYEU0Xk1O7g6DjIYOOLv14csVpezb22eBv/dGkcBLBX4inTuUTe
15tC7BXj4+fchuQ4QuD6knqK+cVWM/H/O8EaY5D0O9WPMy2ExuBJgWnQVz1RHYyDfANLiYQ0fYTc
mt5Otbudyb2MvvXh0rrZURdRPPFPuVMl8cUFjYaFbjRI0CR34xQJsTUZKDkBENSwnEJdDqQib2jp
D+McOCatkoj2HvkSog0iLEoaelEATnIvRgftc3Ov7WA8sKyTpX25Y0pjqgPRr/mwNaTNf1RvSw3a
kvysmi9r5oX0mTGulNw3T0xbUgDssdhZQfsRkE0Ybahb3YlV5Y8+ZXmhsntOT5i7fjPdcMJcIN9s
CiWYgaEbWWkPTZ1SMxUom7lMcpAa6jNsutpzLmXKWspEFHL5noaRdKZYBN76bgitSZ+lkszaJv13
7j4nxHvOiz0q9/NmHOT/xnxHjkqbYzGPzFTUN4HjtUe/4XgQfNexNl0IhBVRNhM9lerH8R9r834B
+7sdzbYSGHm2Dx90bUtCmOqdY2dgk2u1+TGKiWseG9OTN0ezkmoBZJ/9h5IrJ5nMqBMcCOyjnDFL
MIatoGIXCrEKC7pg+DiOI/ReIa2eCbDYrryW/bBUIaznOVw8lQc+gqHZQXlmbD9B6qapXsm5HqD8
8edGAVgiTIukpYvoXE/Eq43EaQm4bYwGh9j4HutQYUupFVs2oLZfCj3QFJ2A+HXLJc+h9ZKhtwcG
p7ZbOniy2UXhcedssCUBiMY7YuZpdceTT7oPHRNIiBJtteMxaN83iUauTbnvrTmiFTlBGQZE2eoT
8vhix5iiPAmudNN2/x3uw/Xj/CWEpwxiB4IV5cIKraO393Ct1sfhm36Rp+UnEEdlOMk6+CMTTrBq
TrexvqgrpkORG+NA48DzhcrcEClH9TWnDAGz5L6puaw/x/1pZ6n42x79RJ+2gEH+PGNUxMeAMjYV
0DyL8FdLYibdSH0PG7U315QMYXGyYSVFmbpVD2gN0WitFNaNtZ2a+IUnZyq+uX5aqgTYF5hXQNET
YbJMoKu8Unk+nOnyMri3WigiLxLTpp3mDV8RrnIvhXfmDE+NW1mPO5k56GIaNd/JJMTWWEBN07S1
XlR+QYZeSpL/QI0sgNXlF6OrpoYS4fLW3UIVAjzvQWUCHDF2QWiF/ycoXVLcRzzTfrOACnvR7qks
HjidcubyrYbnCmCgyPvS4f0lHHtVlCuP5K7pAIQmKnQS6Dl/pQorVYcf2WHUApWxpdmpXTYYfBr8
wM2GdPZ1vE31hqO0YS2jWWVs3plhYCtJKwq5cHHSCAnXVFpFIiyCxBbXc415xhFr/uvCHhuPVJe8
jcBXWLFblFIcNnI6nMCnVLrshXvq1Sm6mgKCr3NTuzzQBuR7pe6haoU0j2XgDjuRDXwCZNPdcvUe
gphFHNkhZrjQ3TdgSDr58CBT3AoLk4n+z84rZE6NJx1o8R3BPm8pOqUBgqEbpn/rIw8L9i8efBsw
BULl27k16lJgFOGEf01XWS4zgOFxr1/xpvdHveYDwcGE8nkcxp0FB2u7WdVikhiFM98AVS42IHzP
6qt38k9oZmmuY5D/3YSnM86ecnNJqOBTebiujkyJIUSqFpTTHxPO7cZEPgltOTMOGZtzLIaH6ive
R8xSdNYEX/r4rct9by9WSCqWBdtbm4yP6nq6Aa6+c4tfP5imHAtFgBdbvZc1DLp/flmgs+xaQrIi
e4F+OJWnXLD1HxQhB6GyHmV/GuG0frjZA9hz+D0c9G510xpscdnPQvAJpf1OkuE6syjK68Anm5jM
gS+2S778VPESZfcN37hp8bqLu1b8CJJhtTk5roWryEO0zyMYeOGnqRyWZAFNUe7RfaKnKpxbRHTL
/XE1DqzJKpFqjg0sGPyNdhJUYIEgqwzoeXYYXCnQQcVt8CyqRnll6XPtRPB4fWO/WGD95MFXduQL
QUxNUmbvpUBoJIIfpG2meXdTno48gpyDn56oJYu7P6YpKyqIXZRxBdne9B6k1ZxrMl0jONAVRQwc
Cx+QkvhEp7YnodHDnXM5sM3Ab5QGxYhmfWnmkMxF8vO9y16K/n7JTLKzIOJofZcUcZdMEYDIwYpX
L95Mx9uc0zsql8sMbZGqYCDJx+XwCvhpzTbENBoDwGZ37YWKbPb3ZNSApnOMAfP6MsUT/5ApXE2a
KIIF2bQHDSYzwMb3zgVwm3bHWtaCDgiYqNI8/bkHbDlcBm+3h+0FQxv2rdRUafsMsFzx8DK+cMj2
meg1AkQSDeZM/4CTX6ZlldJk3eUKWoqTC2wCuxU0ByjLGL8Qhj7WCzpfOByfLepex8smaTz5G6Iw
i1CkNhIwfG0fNLsGkGAcwGFMSheAQ7COkyeDsvC19rDYW4xY+jtuorfavQ5drFypI59oNavXqkb+
bV2nr/5onAd7TiSr4LbdwJ8+ht0NUdw+AgFY0tPJjS7rVaBV7lT6zOeJ5rauYDyycyt4UOjZZO7t
vacLFnrmLE7epgNn6WjCRel8ysCEPkUo2nwxjHnrg3K+LoK/TI7TawpQan5UjTPFmSWQM2+cL25b
3Cni1drwyRe4I3E1oGzvotiK+yIiCDcaJg2bKJS8is2r87As4NnDPT4u2ETPl6t9BFAyQVurh2R5
PVoF8ZHnF/9wRDWIcQ3SGOdqKibX0LjIc1hrS4rxL8OcSHA3Mei/4y/lhcgOSsUmFO3te3Op817q
cKvVS2UoTljUS5/mFo0wFwRtEE/B5tkvYFOVIwoEFFBlkZb2jnLefViPYLV+I0xqe/MJUg3VOAvz
10ftEpuNMrEU21Wd0dm5192ETxgsg7Y9yTApv/IU5tq3MXIyFgULYmw9CYx8V9BkfPPA8V5hrnOO
O5v6w9IiPvon2KdYokGUmOn73cWuaWE4gO5+GXo3JBuTTZknfHYYD+ju8xHfoxgypwF6ScPeFwuP
cPHMy1UDtUQp892b6QEc253HM1J2pcbgv+y0xIS02j69tkrJHx/SD3i4QxWGXd9MLFcVAZc0/oR8
FqAUUXApExqPcTBsXXteGWF/uU99j1Gw7sH/S2N8RUiNvtGWVash5dy+u/60u7TVVmf0CL7TJgjG
6FrHb+rutCbfCL4+/el8NWS3OFvwJVcT6IrxYejtiKYPvrTjD6UWchxvBXRiIkz7PJeBMUroT6GR
LzlFG6qCO4kBPDSe/zTisqEckl0PXaAPoD9fn7XcIlCqe2A4JZdzPFhPYLCofuKK54JwJcf5hfOI
tC7NhJVFdpjgPJhFCtpoV42hWa5vRNlGlubUq9tH73vhxPzMNO5MUrB8GSIGQiHI7ou7tDEGvRcd
KqGRGd9RYhSRoieJyvgVfXIdtYgEe9BgBFsigJ5xZobrGJgtmqmQkGmfXtlxCV3G0a+d7rrcGB2N
N9VO3folM2K/g6yobzN/mtv4gFwFCkT1oKWV2Y6Me/2HY+9VC53kQtxmOMlXzlEetOl4UBrqR8cy
64ah1MyibOl8VB8NMKZw1MgEaXg1wnnkJCt+IUbEkoYWOySeI1tCmdaya+Kp+xFm/5LbqdkGq2NW
JWzV3OOZGDbo+8zDfA3z7/Q6lY4XmC9wysXPMEkEmAXO8DWFKIQ84Cjuxtw9y3NgpqxvH7pVXT6/
2TniB0i2QdQwjmzw7a2aU1l9UigIB4QoU0+sQwJN/Lq2YdPrc1Njcfdyrm4qvToiZIKGtpBji9Gj
Kiabc+jh6voTxW5tlpBgHqdyF3udLnT+zENXCsmBJFvwJyYWmvw9H+Z6UiZyWPe/Yz3/PiuCIJ8f
ismR5l/Wh9jS4N4AGRP43rHMljnjGd2t1FYzbAPJS/oArAazxU8vFbOdUef8k3Qc6QTAw1I1jp3z
XG4q1kDvZBeOL3emZhfVCdd1qPdMLAaU4Aa4/JsOccxcvONKOhQIpSVyj+MDm0P5RYT/T5pKqU4g
RFsIeuHHrLvkPOGmU4OSgDuKpZrE2S1REGKv1YJYVnmQZkDNTcbdR9Ff6wJ31TR0OU69oG88JQCS
lAN8f/llJnx85JfMSdu4J8Kkhl/DKZlLvYPeu8f0aA4rnYYqzgO5IpNxr/cmCm52Rom/7ndjlICP
obXizRXfOOyryN16xXB7KcGRrFbutWKGW/vZxdzDtLh1q8lvJELTsevZD+wknoxLDQXDtT0jhNDy
hyqBqoodKOmlvHWBOm0IffpTvwWBKJqvhbodzrJThQ/PEnudzsi0ZhUWKMDWoEuRS9401ckZ5oKt
Y9bFDn9USwoEFVsW7k3NgULxrbSM4w3qrA8SQl8BFh7swNYe18O/i6LUKoUqV1fJABDmkGmf4MYi
3Nv/e3eT6vO2D56qfmOzGr0vSQnVxLJa3NL/PcRoVLbMqsHFgWHkRm1rh+WYJIhRPtd2ptm1qqjO
WbFSlvYlL8fPcrOqvW8EOt0M/lNsnUx1Mmt84T4HhHpQk+ngK9JUi8YZOl6SFOn/hj7ofemBNfNz
N4iwgqekyf4Y+G+pLNd8TSSGeuQ5HrTMZbKmVTw/qspOlRkjc/qc3o0KcaADkstjHfeBEhaG7nkM
kWkOu/l1CRKVggXTn9srakqv6yRuklktiJbQeM44ktGrru4bSAvn2R9BZ9RhKhc15fvHvvo27kNJ
lPgcm6G1CJOplG7TsJ5EseXt7l03wuLBtI93CqJEwHa22Y3cVX4s5qBVyTcQUgA6DDQc4icHeIW2
IfKv+0SDcsoW88wYBA0NE2D+RGJ9PQRiW5ljWO2E9QACkSI3Pgvd3jBd2o3rtz93XS9N2S+F7n80
GGWhtc4Wv2r2OuenPGtCkucWKah683vyTJt2R/Dudyj6pI0i4NPyoGtgM6cQ4sLw2ri1Axb+WfEM
xPs0m/6IZSaTkEUOLqV8zVv6K9GIepeRzjiKKcjVu0IluW2pxjq14JyhoDoelraLR6Od+JFGck5l
jFMDgYoUTPJGU75WAZMFhubE3AK235UurDBtGomB6U7j0PbfnRrhu5yfxQxt6tye8CP6OyPOfNLE
siFsvm/vpASSgWEK+RdiKy0XFEVRYavqerVAnudPAFYlUpU4LSR8Aq/rWaCsABjU0HYWLLCNbjEb
ukitVd8sfcOtEgJSiyfZUq1i6kQAPrjN7vRRH7j7x3F404XwmSoQiPwAKZu7PpFOBrk72adkK5hC
yj/C7KR9TA9V4g+zOqhsm+mmvQU29jYFFVC7CNmSktcTaljfsRW5To6sZ1JlTDenpZ5ekD8Iz8NM
qoQi4Fa8MkPA8HLyKaaCWs9dpsxtoJ66a94r2CdVpOq98JxDnFLSjamQRbpZ0yHhxztbPdE0ZcsE
L8FE8i0pT3zyVD/x66e+lVReazkBzsl/k9iOmavSVQueWPYAQ3eaaI6kfZqUU1+yCTPf2Tpyyy3w
aOr/YEoPx7p7tPZ9aeQ7T5Fmm0GuFoPu0jHBsLWJd3YeHXbxehqt5ezOD+yrRTJ6+H53Cs8GohAS
wjI5yW7PihKy4mHyC0UsvKq+gt3GnQMfNZJprB68PFWTTHgrX7xr3wWtcPXd/TSTjL+/u9EJPGhE
/MjVOlxjVnis5Ns3TMTjDeTC9ovj0AyafJnuNcAB88p0RTes1PyM3IBInDIaMYAnkr+QipBpEWOP
GFSLm9pYpkj4DvaGfPnnlZAIq441qSCh9qJ7uSpyF+yeMwKxJhSo+2wvUFYBMwC8hpjL3LIoM8G1
BfOgju4XtXcle2G5ufjlSk8F235ApKrl9jev32PjnU9ymZtwiTwQnaERNnLifK9ohuS96+uMjtXc
Jb8vB9Bxzjicq0SpkWhizDgPlWCf+354nPSQyxd7T7qREFUfSZM0ZY1jBdv1LLBTS3QGervf0agt
nBQBI/lyiKvqRFzYeT4LLQuBHPWSOLKeqaW+Vqo3mSWM3YkTi8/NdZCkd4MOBc6kQ6q19nJByon+
Vdvv72SUJALbMB9+853DkqNIJ6SeWvNWlIrwQ2r4OOamR3FwAL/9DyeTA2e6CayZXV5EiEh1W0+m
HZIR1Ww26v0eGaOb9X+cTCt7WHsgvOc1k7ET9Hx/3lPb6XCQknRXyD5R34xzSmYhrk7MPrbYzkm3
HTI8pN8n8BkAnSDpUEDu+NO0fPebjDGsCSfaTyC6O4sEnF3V19fxlHKVFpfP7kOY5n6ZK0g5pR3V
R4ceuDd9H9RksdENd+QrFqgaKr9C6eivKH0CfFBwzxp3GVzzzriiV5jYWXVGdi/yQlHI1Vl3YbJy
RKbL68uFh3G7upi6M0gUQqFVg43dCSmrPVwrzrHWOtHVOLHOC8kh4iqrLZcVjuVdNjlMgIeuOZaU
o4UoW5S/iudqbtdgoPogrhQMuESBi7kUt2+6yuLW4qtXCx3wAgCYxQqqRlEi8LayvIFEmzkHybvE
WDkFyR0hmFibeS0fRdqOC6GrMCkHuVRkAsd/YNjVpJ/Hkr7hn/Y9XnU7HuGx01doeLD4/Q4tGdWZ
9ds0dECQ8BoQuRFY2sjJHHwQkXZC6YV+2oIVebSgOJrJd5yeWVOdrf0Ow1VPuYs0kb09oLnFiEzm
+YypoO0CmsEE1podX+AVCCBbUvtbywkxiN3m4nMLDVvgF62vvfzLojdZUEBZuAXtFVXADVSi3fcd
2yngsYucZVwkSi72UT1E9iZ15Yu2iP2XOrnk/EwUUfPOhmSkQFqyCwoKb66xJDvcx8+v2BEmxxFZ
LKtGPhxtsM/ge35vjdQrmzuDtwkDAESoNNSbtVTMmoi2a3lFSGFsb7v9Iqaen2T8yjgXNzxnxVku
qWMWaUARh3GoCXXONQh+KCCrejNS2hc2STLDMPtvGCKs7200hSdJgg1R8OYhgfBLvCiOI2baIWGe
9UsYLTh6KxSQcxdYiiUXppAQfkS3dZ8nwOD7sxqTfwmo34k7y6DEzZ+WfSnhTGUPbVmkQLbxOFs/
YkhBidO+vCiAmt49ypUlbrmVT44AaVpCVpWUW1tl2NynasO1p9DxBL3hB///gl4aGBgGqqy3lrvM
Zw5q4mMpg/DZo9VvewxZPa4JcfOfNj2LFfsUe0BaL2k8tpUF/WTGoj9ACBGVIv1oTxPA5n2+CAAP
eM4b6awXcAMUJTmbryg6gWKv7u+qYoNf1mP3Ie9fEnyzunJRRPmWdZsop+cOkHI4Gub6QJTVStwS
fGBYD7w8hnR6t6EUeOdCW/ZCWh9RcFE/UQ9kyw17JGHO1ietGM24NFGo6toa42LVoLqWQufL1KMP
/WgS5UQkSgVIbqUxIHjdnYNADb9rGIA/NMUTe4VUGGw1gwrZ5+1p/+es3X6DOrFMs+XscAsc6Cs8
sy7mDMuiu/1Xq4b2BWu4RAuuOHEpEFFrbWBfJBzofXR9GrFtiS/nGq0pI/a20pXqc+U9A8X6FqCJ
3tdw+8p0dgcyvTh09hnX73TzHKPbqHRoUCIR4Dv7oqtQD159eqsqYRl7QnqyMSABI4y04ajpYHeq
U3ECiY8QIQOVCqyLl/u9D9bWPo+XOFfYvWHJmJaZgid7Zci2SSgtpVIrj8yGBhDO5S/o6BLfwdD1
1rMcqFJSkQSMjgowkPj7Z/4n9agnrgn+pPFG3/U6bZdDlPIIr5T/z7qncWXvJMWs4mzzAd2uoykK
LynphYJ+8pP5+BKTm0ve917ZBKAUYms71wDgdTzXRmG/JpE2Snrf1BmfwFAFqiqwKz4juT43VdbH
jCQt9HdhsCvelC6ekAmqAQYjgS4O1y45MJTRjXnRjTnaCljyMI0eoJQtkYdPi0sE/MW5z5ca9YdK
O3srfDyyitGLcUh93h5cffbG3fvMK3wexW4WiTKeWXKrdf1+LkSqcYrbXqVjmyEIiwsnG3yA++Uf
5XR0CYkr5ipQ6niGMX7zhSwlyKPbN2gY9+s6o85E3fXf5tRAhvBRJkfk25VsvG0zbr0DwNujzAWf
x9HC5IRTAAo1xST+/j51wa8/e8furfYI0Fhr76oqkgHS9NAs50mrVScsoEU/9NgxI3seBJNvbUUX
DvsaMTlp1dyJLPEDNHFfn+SqLB6BnUZhEuOvDVeqPeAGEKALVpTgeb6pR9Ra5+lOxfbWL8gTJQvC
miLqajIpncmxsXix8mTtsSaCZpmWBfzNFpDi9kX1upEr0hCpmOXwVNB00A2zSnfEiACW2E9AQg5q
dz1qdqd2chUdncWByV14wNGkucped1LHf70KjM2c7FSbq7OTjLuntcRXqbKgG31Zo/RJ/PM47v1u
QuJvGYu7iyCFQm9/iIy5EUJdsc33j5R92zR8FXDGAylVXshpCsO31KSa4TnKg5d9/bHeT4eIkx1v
gN3Vq7GxyvHm0w+icRTDrQV3zM+mYwRqtP5UnBoiStfM1f5p7I+9xNesnkbgDYOIFbqstZgqjekX
tMEDPkOw3hN9/pLB0mKYHVrAdzdySSodkX/B6KMm0WKO4xvvByjdDx2sloiIQP1R4+mxfcqJFXgZ
OPe4PIDbmKy2bgyITBAZJC3tYqWg0kqmWoMb/xgU62eXi82bFAn+cbmCfk4jGojzb5JpgdWI36bx
pgO2i9KiLaLoqdeVwLjsTcIvF1HtlCGE9/1FQJ63BaYvZlvbXSYnhwWlxPwFAxUp/iMw4JZYwgLc
gTObRjmwC3mfhdXq8OYQLuKuX9JVnt8p+u2+fxZjSlCzz5D63tZw6zEkDb7zR5slfXv27NUEOPpQ
ylrQeQi7LOwFmPB2FA5JGpdVpw8pHgJbtT98dczsZCkLxOgpehTHaHdh2D5Me91Khk/A7/fACHSx
wakoxkLC7RQcLJ36pBcznFYrGkSt8zxIqVPXmK0xtu9PJ1lIU8hJdPV5+B7NSX7/FfYtrPS1hLuN
m2WgIpO7EKM+UbXfWOAYlQkR1jB9mrUg2SM3gRheBitsOtGvnXo8kbR3Tiye3/XrtEqHxKSMakCC
UjeDg0htMIDK8CwDZAyUBSXz+c7w6f9PcpDoUoehkG5VnCJYcfLJc3XYLMws1PKuUURqMdKncL1E
5Dw/Ld/vcAObcmlMURArCSOrpT4zwLDN8A1Uxn9AfWRYyPoUKp2gosUT2BK2TzCrpnMZsiGhBa9H
SEcZ5SjMysUFUSSX1wY29eBb/CrTVlwAgpoL6ioD4a58JnndgtV3lAUA9KezGNcRCp/bHJTAzMth
zskBVBFl8wSgqfEIsdZJvej/5OMyz91ABOWof/tiEZj8f7WRQhIbzsVbeac1QTu05bVChDqNjcWp
IBCaegC6jq+g7fRHoVPGhR9pscVQz1+4b6tsjpjjsEF1Hzy8uSpGiUnm/s0tLyCDK7YatTz1uoFb
zRvSfM7XB0dgXTRcI0eUAA11GK2iI8OkxjaWK1cy5WMXOuMyKukr9OUl5ntqIjFVcSXmeo2Qoknr
L0ibRWF60JPjza1+JQ52Q8W0CiPVddyvn49TFKwQnIVjNvV/a8lTGQS3+PiZgCjZf6bj2SUmTrBV
WReB65rgojuMNru2pK2CiCJz06fHwreO8HK9iqG8/CGsIjCjelrxayfuxOl48ztzTaKLbpAH8CPp
rJkTaonFZTOLHj67WXdlfCh49M7OB+nozXiVYhO73O/zargsewgEhYGj7XOUAHzW5cB6vNkKH5/O
AckhYJZqOGXXrVAIatI3fplq1q0P91ZMbl+Xwyi3T1zWf8T254GVY1/WdsTROYo+73QfustDyVCt
UZXUSAgvKF+4o59c3blg5Mb3LxK++0uyoiHATZq3llOP8ly78YMqnKNtRtJrQ44EDb7Y+wWNiyrx
GhsukEf8Fm+rT+ZU8jHKkNLTuXfCWwLd0j+tB6ajOpOB5/gj7wtOyJIJGIU4AAITsVBT9ZQauzNl
aqIxH1H5c1ZWBF70UdVrLgBZCIP5F6XeUDPMRHJa0fG5viCzb5cwNH68dapplgBln+2jXuxC3W7o
+rwOHuDCnsbEUlnT6K/2S3gvtIIFfx2iZ6DQKMr+ohkZuguKrspyaAd4GfZ3zNYkeV4vpuN2YQr4
Zem7TU6C4A2Fb6BaY570JrFEXCFo9GnDpBRUR78mhK8MXiG7DyHsshDgG1srHjl530zFQqJj3xSj
swH0O6tdGuGjwHZbagV9gjOZBCW0TngeiP9pMe8DppdGIbQnQB23syFLa9plkM/jTwEH9ssrndAH
E/HJRIfOtJMWUrzpcjPMYI5ShpLXw0gc8k/6C97Y/BFf+ye7XCHfKQnWHBydclS0KnChNX9+Y6ow
dMDRR3tSoITWVlIT10v+6w1lzkLiL4DPV1cffGtMV8tifd9PS5ORJlTZ2tr6pmhm3yMTHEdk/PkJ
t5mqOOFttdzHhfFKcJUOG6x+gwKSfnQ+/ndq05k42ZTByPIm2IU550RIGNJbkvS1y0ZFn8ohBmEg
4/5fg09AFZ9cFYNogmcK9AuSQ0eJt+lC+aw1Wy5vCZwCVI4iRmDJnN5G99rdzGm4ML34yYzVq/SY
S4ma8PdNYRCZpHB2XR+FxWqg2sghcmfh/vH+i+/vb8KC5sFHnt4Yqjw3Y75e794hbx3D+9HnA8Bo
uDypr75elQj8HC5sFj3BlJGQoeg6EYoCV7I7koHDaVHGftb+VPwiX4vE2a3oNuof7F1glskzayxS
xkI6RO3p0QB711carViYAD7ifzBFF1USNdjXZz3Wp6P4+Ico0HqYy0I9b8rx7lJlzxil/wert7C+
B0Q6aVAJqqee4B7YIJ9chYoeiBy6judqLHxzapIhPzl0NzT/5Ac693YpoXA/0o0Ukqt34HFN2Kui
9gnGom64C9395WAKfWd35EVFNEOlnLcVAg+ostRZAL3opbGLIzLT2JCftczxgr4oGNu7k7yhbkJ4
s+xllZvEVt2HRlaTzj3A9vSc5j0Wg/EhmcV+1EvP1S2M9vR+T9nv5WzJauajhvy31NGz/eQH5cXV
hGwg/a3FO90GmGjoESNLPfc0NAx91Eng6Wn3q72yMZvbZ7K6+qbGvYXyrknjx5WmrpO/CZGGemYr
X/qWeUU5B3eb7gYF511iE7DxrameCKwFFrDnLTiVMjoFyRADzOoAKe8VSnLSq13zXK3VUAQaQE1i
5Ucxcx8amAUbTQ7jqcaTaPuHrICWzm8VyxbbBsSK1b4rMm9nK1xbfM3YRC577KDAB6gK0gsULZcL
tlwCssG/AyuV/KW+L8rM7xlMjUKldTtqriyBIVa7X+C0rhDe6UQyy7iJrPdut79PpMeJbJGrijxQ
nCzaADVtZv9yxRseiaxRM111pc/q/XHkzRMgyeA/H5tSCubTjPuZQKjvO8zbkC6DDXE0yZ5TSEe4
qaPlJGPOfJiFLVvprnLyXjeDwF8oY5QkfIWIP8Ly6sGZMOkOJIzKK96Ns9sl5UvFAA1cDn7ZLKBT
d7qOFceeusUIMdxRi91Zwyhf+SLpyeW65rb2mZGEYMBR97VOzehLGWFlIVi5Qxh0WCaxCrGJ53s+
leqmS787Xpg6T53b4Q114MyZjWkPrtCbJZ61TYlVeKyG/om2JX5/adTcyKciUOMJPm7C7SxTWEqo
8OPpy4pmmoN8LRm/pfkdreRsxEKJ/gG9HmZwIQ7zFlhEbqJBkpaGMyN/iQKlThtx+6b8ptmD4W+g
C8M3FMc1T5dNRfftTIaRVze2T+qBmI4TEevLCyPo3CPgVh8tW0o6CMjvh3KCAqhbMP+DeXpXQeoJ
E96yWxndlkYMz6lUL4KifbQ7pToLM3rlWXawRS18jJSKnj0pg4sf1+8v/iaAVUWQhCofadlNHdlk
qU3JrlcCdWsC24cNgZfhB+vaL1RtWDe7ddkPLt2dPiZjiDkb8VOOv4gMAeM/kMvfnKktVxZ016Xt
RRaYYzwrdC4eOvBPiRtlOG6ifdROapv7T3/YXcyJ26eUg6QGTJAmFuPXD0sWOk6p4ALQwbkpo80h
/4rgVNlsL9ZOW5kLR1OZ68iI2KP+5mvMsgkQSINNgCbSTOf52CML1/jpYCpnRbY37kXzFClSCdNr
wvANW1D4Lm0xrvvs6nw7qo2/lOD+AVaVCV5rxAxbAzvGlyyk6IzNxaSg7qOCDZW16WSAIwM0gYCS
ncHfAEyfiuVQtuv5XZdOBdwA78t65jVT/BinRd+oa2XvNddVhDtmuit+llum1E2sH0yehAms+PEA
Wjlf2CxZx95lMWAjFBRrUfWcDCj4h1jZPcF2PNEW5Nnm9Ip8I5faLkG/0H/ddZc8iMslH27ZeLsi
EYxoZPZhp+cDFBtgxoh9JtnveLBm1Ovh900LjKa9ePzVjlgQY/ahmENEHCcPv0Nhee2N2WPDcyoM
Gy4aimiUaurqLo6Z+1ptmsznaBnHmPqnyI7RI2GohYNI8h7AhFk+ezPGBSOvQjvpbXA+QTCE9H9D
t2DxxC0OKKczH7aF3zw7a6Zc5CIg7VdefULKW7AF1eLgGabliJqY7ZNZ6x2LKQ/3AgbwotnNjuJA
ICWbI1pNom4LEpjoB+PtDKj3lpRKdMx39uoZKl7xSUMHrlPM0Uj5AjcoAjzFGbHvFf30dSRawysc
Bc86YYgvedsyQC2sH34gMXel21oHtS3m0pkfqaV1D9JuTtpLOHJwkKGP3XcoHnD74c+cYihR4gbv
nI5BD9UP9bgqSuSFaNaQ0E34p+Pbs9SHAX0Tfx5AFQ3lVp0FOkz369jzpFizKBDE0Gd18A2NObU7
eSylMSCiM8hstAofRpoOA3kID8BZvP19Em9fWBuND+8SCrukklc5P1Y9T/qOKVqCxfWjmtt0k7MF
x5byX/X/C3BzPK+IKARAbV2imldyGvpPHWJj6m0Y0kFsNFoCeCFetG+UiC7dq9CLhUYCBmx5aqa7
fXzG5eRHhYCVLOXFK8W8AIgD83dJDbwrM63tWKMKXfzVvOuqmWkMKByZjXNESVHIzFNjivm4vYfi
SK7XtQEHqcLuwSdSKH3vWiZ1XyI5Xa5KZelpP1SvNxWhFzkkDmwjCDyKKOVH6RHyp/BJSnExX+NQ
eIg881q8EA68nVixjejogRdfv1AUCbV6wKAAlW7pr7C0p/N3m8LOMasmuJNsxNJtlAdtnW1iWnUy
fvMZ7tXfvCNiTGVzeQijPzfPadDje7Ox+wPfXZWGsBfNDrJdqUXdq3DupaTX5OP/4tI5MjoRuTiX
TTPDm0RMAR/6XeO0CVbnO13VlQhxOtM9qYAB/wtKWgYHv23szLSvByxEfjhC7xFzd6053bhq6VL0
dCNYt9HWeUXVBhUzknnGWwrEPL1XFSoDc+KxGQZQlFROBmRN3pbrfMh7pJNHY9DEdMYA7BzANasx
0tSb+j5t0NxEQXA/I0dsTRtATgZu2aZNjkJ7AsbNRCEWlvdX8KClphOiGRcWo28ESjSoFFlHbaNL
XgjlV/MR6XCtia4IhcF/RLehApx8INOZ5S41j26xS+28UR+zRH6XIqGxxzIloxvhHr4AscWKF2VB
GaHcoNqun/YYlufw1iKWsOqw29OJIiPTyCdlWCi+yhSiwQAHSHpIotNeu2PzuPHu0zenJW/l2bg7
UQ/Q7uoJQRtbzlS7jAhAcxLAz4l3bEygibpC2S76SjDcf8QrxEEpQ78vJ8tCXkTnLnr6F7RFPiEi
FnBLFt72Gek1xwQyVVkYdil+fEnfYJSQ+HSf0ge7ADc7ygexRhCSQM2UdisA2UR3PgBbMEyATV0X
j7kYOtWyMG+aj3FCQU5DnBIMQSQQfBPAqr9Ww56A+9INMPkNfQ5/eu0WTxDbO7h9l4bSVX+MV69n
J9OHA9HK4K9Y+g8pJFVV+GY1RCxnVqNmO+a3RpENqFCLoYHRnSnBvhxWDRwopjQH8AC/lkhV9VRO
ZO9DMwT01XwoNmoCUtLNVkqn5WsubjNx1BzeBvchaw//wF9mrLn56C+WNb2j+BO2jawQlQIKeLWv
F8pSHvQky87fiiIv/esM2M7Xa9at9qOY+lQZd3qZpslm0UcmpgbeufLgAY+Q4XUMUsMpFL5QPlDi
TztJsKBu2KFi9WhAbU4RKGUP6pXhSdZOVc4SEkyK5M+8BnY4MpNDAxXbkSXsm2F7uE9b0MdKVvdN
UBqrD9qmNjYZgKfnCZ6Nfznb+dvaxtpdUqGEJ5EFwViBtyEmAOI3A4wxgJ3yNph3s25ksFnC0QZX
xpxN47/Qb68/M/iXpgzR0E6zZzZGRWEfjskpNLf0EicEegua9kZ0VcLHGgRNxocx9Wqj9bSD23Aj
+IMFXPBzPQRIRzja9q5p4uJfNEKr1t/p38jUPdJOT1IFSnzjZqYseDAAcLYYb/zZ1y9+5kSBPfqx
MOLA1Al4IgS8s91FGzJOpCnVYj1L2N1odLc+EbYnfweif0mjmPTyTw5UhQLEee0nRnguEw0kAYvy
3I/L8OuB8Lw3IHch7RixsG6jpfO7awsFQlAr6Qp+in9/0Ciwl1c2HItPfT7vvbynVzEc3ULgJ7zY
+roGioAqXhvqXXKmPD3fzXHk0Hlvucq3NY5j9qHdiijUIZ9f8sWgThRC39aGo8KcKtR//pJgSxw6
FzDRtgOqZl4P30P6zfLMAwEKTm3wP9iNU1IKqf6cp7/qen/d/ot9RPDG4+UYHuyTpLm+19GBjmak
CtMu+2AN9+mzaSzRv8uaOclvmdmeNXGrw0+WLuX4WGf/9mZ7GQzvcttiq6/gyCCN1yg3wUgAA2pa
x3aeCG5nKQ3X53DcnkI890JMCdZbCYIepi++fZstc1k5V9R0JaFA51uwZ+8S7MqRGQ4zzojr/idf
isOA0m+1uH03ZVs8KqmdtOU+zLQ/fxGWxgUmNYbbgY0BeGb8g4xkunP2m4hZv7UE4GzsQJ439Zrz
HNKnrsqGmMU/A4yScG8hpUa1xnYmZuQrJOLaCm1NfADPBYZGxxeSrJCgWET5yaT2lAOGG4tvAfxS
1EjGM7+7Ke54lUOUb7IdVqs1/nkISfCX9Xyx0K35dvs2YfJfXfVcoJn2TILSldGxho/z32CD+w5T
p/WzOF7jWdY+Ixl8WLEtRxJ3X/W61U2Ppl+nJqIIRISB5Rqf1txXQ/0BWQBNLkrES0D0sMR762+O
F/bWUqc+TEa+RKYzekmIrBn8J/09ZhOyIzahRhyBRWoW98PeQWEIW+qGYjnSi/OMl/eT1z9AYSPR
SOezpdRpW7t4ZWpyfORRXsGK2oO1UtGyVXCWFhoFTpq56ECchQrqte88M+OdmYhlfrT5RRVpuwDd
uiQEHdXLpqisss9AcudmhT5xy+35iZrSIWeTdWORHwam4b8CmM8gF8KoS9ndDPTEAIybw5mDjaaB
wQORe4oH+65gAUmUEQmi/iAzQ4CP7C6Cuzltp9pVH9CKiENGEkto2Dpv9+PoGcteg0250M+CxiXL
WEQiz/XoAQxkJmQT5b/khTMdYp9Gj/S3/56fmIEwgS8s/jVJPaUed8fEDHwD7U2h4pI5+yiw31Fr
gAgGSHOiSRawGjnj0o4ehSpUz7rhTRdHDbo2vtccwcreG7djediFpGjpQLDjuXGR2CBzVZHnwwou
FphYmxkqBqqdvfvAU2ecBu48HFjYS0U+zLtJHHhOQOfW6et8zRfZZwPD6UNVIVAMbc8vKjf2i3qL
luZ3e+14H/iNJ67NqZ/Wv75zpDlrjll7SbmLL/4AkYGkl71qgqDiYS166//SvvyckjaGGu6lAJXw
dMph7XnWCw9cGohyXitumjuot8q+QMZg63SsHD8WWvjZr0Fzg9If+HS7kXWt2/BrP64F8smXCEOe
2ROkxWNmZEtLz1ojl/rQTLlvOWVH1lIQ/fILXC9/HSFiHSeOcUWnXd3JEbPFYeFVbir0fokyqS3n
gAhI42wWcpbGXkXJleziRylrdYV2ftGjiwszBxnjnG5fq4nr74/9RxR4MczyN4aF6EmlOrwqse/T
Cp9LslRymvZqGGeywVZlM4vh2ayGqHg1Y9IIkdOdb8bnX9DZxMkZaZ09Gmg5ADYdxcsYdXUB60iy
S2LOjBs9xRyfisBnuCmlekwHYb++53bBB1zoWfq3vw5PY9VHsARTK14IPAvJ9ikUuVpHY3cJwP+M
DdPmvSwYhM5KOewulXoQNe/vtm8UlkpM38y2bcIUY+mohNDLHI7zmJLRvFyleEMZuP/HdMMTc5+g
fOTtBbuYytMhbs9JLAIX/0b4ULyw+yqpuadElWdHDmQU8vnE7ccpjJYbpB7413ufkxWjjqfI8zwX
yWxvDyIHZdeJxdglRdy/hekTEMleDWNCi3+XN7IR57aF3G4SFNQ5XcXmozzJoe6EYFNW4zjb/aFt
Fhs7ePzGJTCr/BY04qKp8Z+S5eJj21iVATJ+CQxJJJYmyJioqghHSzvJQYxbX6S/FFtF0XK6rUA/
RwCLgsB3yPJh0ZGq7/K2iSxTUdr0PNbqwqk53/JZlnC7aZQx0wXTAmvOwHVe23/jI84KJLdNNU7p
tj6KU6bjhgGh5voZjCPxOti04b7BEgmRxlx5NdGgbaFXaOhfKUR3s++s9c3rD5SFvN89IBMHJ7ac
L7tVu/EOztUsYPqeOF9AHmJRjPGNqTnV4ZxbeMFgQabieEhjh8FMSyET6Lo1cd2/nm7peb8rWbNE
uELYTjTbQc+9uoWgwsuf3ggkbo2xo49EZMIGMkElpqk8+0Pr4hEuxAX8SF3i+zon0TGr1Isc1R0P
YBuq+6L5Y0IywutR+zzOAt3TABc0GgMqU+RxpnqNLRtd/cUZZNFw6B2+3hSQnUK5e+EeJLEQTcH7
TrJFJV2MguPd7Z/AGrlZNSk88Ke9CpkOnxvIxlP7MiNeWPN7JTXpkMtejejSCS1kiwyvOy256u+t
chzJOYCysdKByOujHBbAwMIRENFIh32Ysc6L3xzZaZtPQ/2T13LFHRJkZN7TERJEEZo1rF3XeM0G
+vaVy0a2HzN7SGBuWcwi2C5U7W05lLcjnuBXEL6iRiyIp5nKeOGJgHp8k5NpoTSGhpeD98a8/pgi
GgEiDd8JYksMWsC+g2a6UANATiL06i+p8P1yb0dG4VizxAzhnoDkLI824Ig3VOaRxV0fbXNqRvUF
aqzJI7Hj6OguJj3gWQ6xOVqsjCeX94hj6qB7KKIXHkm6JVkbly5LIQDgB7UUjRqjSlU2qSC5NJFB
T88fBozynszCgq61a30zBozS1U3M/dY2jaBdjAJoABDgF7TdQwR3bOf6yVpIj8QroCEGOAhQv5TT
l3/TNwNDO8aksMHfoe4NWKw2L6OEgkVSZIMlXxAo+YP/SiUbKnUkqARG5Fz3ppJhBPdz8gqWOtT/
tpTD2J5DttKkqh5aNYZn9xp/vQI57Q6cFjcSbgiDCIYbkr+3kIGDjiPf/HEZQuAKJs6MdRciY6PT
ZliEmxM5KQqYS/Z8mYVZ9OwUKvU2JRl4xZLfLSrASo0rP8+feYkIv92lduFSy9FqBtegJCx9CL2C
wleEgA8z/JKtndVztWlrY+OGyH59DvsMiGpKm6BTPP3A7GG3CUI6Mym8IR2nJ5ogXtFF/U3n19eR
fu/K+V7/d1AKh9lkPAEtabHJkDY6U4862tZvqPLgLSGBba5zQ416gZWY7pZBm3B9QFshy+VC+7mO
3k57VCsYxG6R+SkMY6+k0pT9aE068VswYdpObQldu3jOsi68Io0jewIj/LKABQsWwEan4WSouVtv
GX0J+OKWdWSOhKZvqP7bME+/FDqDbn3JE0t8EnPVUb2+8mocwhj8g869dM9STfwoNS2GjIUcRGSr
6vqxSFqW3aM3sADQIaQ5+uExy+HJVWNgcFSQOZx1xixS9xLsgZVIjAhD1jVBy9Jr4pjiOqgsKCDC
4vKFLn0G5kG+yqkDD7Y/QU23mGq1YkBxAq0UHCLDcVy75RAX9ilUrfES5NAbig26M23j3Rq+Ep1n
mvM5+dDBQFxrSZPVYYI8drsJOgW2W59KyqyD3VwswLifzoFC2viCrq2kipWcDYKM/XCPlVbePe6G
rRcibhdg/Tjz6H+/FFG1fv1AhaFO2bXcArf1YGU1MUQwV+UQzN88TUB4g8tYDmX3oqPm1kvEWR7F
JoMgWx/+zR6J8Xy15iD6JY83WOg80cev5/Vy22X8QWGUwp7lv/dmPrQdnEIbfWFkv7H+4p7RQsdp
8vbqIrWXCR+HueZd6R7Q+PxMLYETCIkrIo+PNmW2Mc9gH8S0/7v0PD8ar2pWzMo9a93OQaNsPtDK
85o1CmnXKqgA59NvyZRDHY+e5EWQZv19zZU+nCh29ujHPGa+Y3hPVhw0s0TM0DN8REdShQy/ILp5
62Ws+nzA7T9Vbts/bJkZ1pUxBRjVykMLCKalQuqELD4qk3hBS6XIet3TEMHQns+z907wElBXWp7N
BXtN3e79k6VkRBo0hqK5NBeJxA4zyoKd6KMb0Lt1oxXuhSp7LvDaZmi3kfistVKzZ/3Qb0CRV/Zp
U6Ik6aJNOH28vWOYBDxCiZFYspt0ZWFWj1WywDfft3DgJSEOdQrLab7Z3pbuj19I9yRt07XBp72b
ApqWG6XUuKsu3wMmAo4HCCkt8O1gZNh+VP+Dw6JMPdORkgXY/hMaS2jxmnQwcQUaJicHgbmE9OEN
ZN1lGYwHFe16DELB6uAlFScfaE717BVXGCrJVBbmXucKviqo1nIsVwo1TPuZ8EiM3qpYzcyQ4UTQ
VLnJRw0gjP2q/MURIPTUE0psryCqJ9QzZyXV01exP/5h8OmtL81Gr7ZGycvMIzQh3Q/tD/+Rvb7B
HkhM/sLKdWCw1QO3Wlx4NGMvMv1XbHTd+cgMivyOOHcCi+K/D4YW6iv/Z+5W6MqOUv78symP450m
ux4bOg+a0k9S8ZbWsuBpNLGEfxsURUIl6buAJlrG35CWhVa3XpC8bKmJcS4reFieiOvQKY0yvObV
8rgFkTaSycFtEQCghz9lKfoC9gRBLIacm5OS+m1vc+MbDdT5Z2aY1Pqkm/c1hrGLGm2rVr++0h+L
uBDiIw8b4i2c6a+YuEbSj8bnui2R+RAx6dWcPiKpx9EQQfIngzbxgw8BzOCQd8s+MAsWikkbVdir
DKtSC584k+YeQnamSd0pje8sK0N8p5TfppEd1J2WoSfDpR5Ey6CmaoK9bPW8EtAS0koNHK5MEJrD
IFil1RW1u2MDNQcDWEWnK1hJB7ArTHzs/hdJa5LCjp7dJutQhVYQ7niPr6dq1kLWRUauE4O/H+IS
xnXAiwMBC99CRf4uqecZmmYa4ZXOF47OXqTTEADNtibQW40IWV2LMEK9qlcjq7Q/WZtTsu9wWxG4
ET4jBGbCKZxR0rrt9BkD7ejqVLlI6/4YuhETHKZM1ll93R2WmuaiaC3vDq0PzRHVVX8TGp3Ih8KY
xPWvDmJK6YaECjyDbpYZBCFAZ/9zhD4zuXIY6Yzf1zA1B/M9erTON+KTQBo9NKbiNPtjld6Tt4+l
zJFZrETpS6GzEAHeLTqN17fxWmJFEGL2gjBPV1eruvligpHGOIGl+4Wqpveu5Ud9m4xQ8FnLq1jd
7o1cteEzdVSbL4SwmeRIgMq5hvbwyJLHi/e5NZ7JwSZnLYn3zGKmCYNmbxYuIis6gbn/4EFQrRxY
pvgkryV9dMkVOgAetQNXVFqGpmSC+gfJowK2ITMD2lmsGRCjUcrug6LiqR0Fk1WNEbWKlr6WkJGx
sYwC9MV/+Sp1vhwcRI+Key50peRIIt44CX1Nxf48+YJR+8+KFCyngPmZg9QDhjl74o14cz7M+olY
nQlTJSdPISPQE32K6xvp28xkjuu1KAEELIYaNviVcZs/dncu0otgJ9OcppEFoYY/s6YGYl0LYbMK
q7jrXEfFoXJLsAVHnSoZNIUtpGUMCZ7Rnnr666USW/pL5/PNoWhZNt/iqi8aEy5oFfvgmYLksxB2
HdotXi8w+z3GFrWK9XlwviFFaZSYTgBTCNcJFzZPUONFPKRedvcL/+gquncAxzvBdZAy4BtzPM1g
mlyyV3tpvSj4OMgLM9/uTxPsLBZKM3IcrMvPe/keqF3MrQ2iLuuyFY/VJQSQSKhBCzy9YiOA0rLv
bmB5qXjfrWz6H0yiK1xqiMOcP8Dv+tTzArhpl3TJIYugfvUfX14CawN415VSxilLvdZrueR7JExQ
v/fJAIYly6yfr3YxbxLGwaoYEY1eQDaKQpY91grib6DCNttVeij9baGkkOKIVqyuHF/lTKt1ML8W
pgEHPSvIGGfIWn4Zb6bVKFvTsi3J2px0vFRS0Sx01M2RT3wUzZdP25aezXR1jXdJR3o59481++1c
w2ov7CYVXLGSjpdqMBxI9lZ1rHiSoO29st1jar2VENTXOCf6fvQw2PBCafVcguSJR8Fs4JUvwEEl
Hg8M+Qw7Acsx7F2GkiH4q2FKr6zMWl6VRrbvN3t7CeiyuMNj6DcUdQnr+yVfzyl37H1XQKpl7utw
H/MfqVXAy9gwitTYr96pe4f9J5ra6Oz/fSERInp4zbuRzI15Co92ijb4sbud3ZrEZh736w230BFF
jojI+CyKdf3eSRrqC8I4EUj/glVNT/uqnTEsY01xbTqtjaTZ1g6mRuI6OZsyj9QZIwbbRnqIZ6xV
iN1Y/H6afnpuvwXu4Jj7CacirroKyGasago7HBFzHxrGnFdG2FeiVdWesEU6gUF8/p7o7zt4is3H
5K7Nlrql2mLjfzIwX0nqaZyDStwB+4V2kQgYjxNeM842VTD7R7RxgZh+XpVt/dQ1EMueISb3aB33
ALIdGENwfIjvUx76SG5hFiu05DcFdmJcT85xKPyosPKdwR38hgmly5o6CdZ0V0fARZryWF9vWiyt
NygoTbx9XRRnuPgjkfJ8y89W7RSn1s0nz7cj/pzu+N9VAN9wc2Tevg4Q29c4UoSGQfeIqhbozFco
f4KTpfNzFz8N4cq20V1UyHtLPVt9xqzkPWagjw2vtZOY2CGF4Zj/NHvdxRMTsNCCMInYwEc8sQaD
81thdALy7xCntBxqujKriuDW2/j3g9pbd2CVo3qGqCaI4QrFrKrbr3+mJv/bJ09eMB3Tl7KvFTOk
XQIET2sirvkoKAahuZYBmScu97+UoGNdRnan4Hn0bkzS/FAPiSmjcBJ8348EZl2/QxNHMTzi8kUF
cnx/dNWUFhz856uiILGN/y0JcAeHYV/UTbes+xFSmVUw3ZdpXG7aXOCQ9IKRQTSErUjPlA68AyKf
5YSQtyPmcdHY0MNiTvHZR1k7fZLFlXLUf8gGgkrLu4GTjgStvsJQseLEMMgcHjU420J+EQEZ+PhP
2VW3C9WugADQzK3aJFU8XzgprbZT5iW2vfC7KJMnNTA2yqHTNZNLCPykRydEuoWl5wkXyyg41cco
uN+1Ldn9l6vWR3Udp5+0y3TiLnUFQC6msdo/oZjsHmr+A0wrTFsKvCeLnvIVCnh49Bh0Yl/nAT0x
3Z/0FKhkXAIf+t96ijolDGuIpOWdzjj0UxaENySA7tEIbJDRGVZdYIGPmTzRP+tF2jcHU0LKQ/M1
gu4eN2efl35XBUO1+IpzCM5iWFI0j3fA6m+DGS+A1ZD5MpKow4d/VDcUWjHcW1wQYgJ3xJKdV9B8
ZpsaqpXydeTPN+3bH7NjkhHNHAc1ifi8HBWHv/FksZwnBAUG4A4nN6UQgBMFwl0YJS6ZEezHhl6V
trUZGDVBRzqc7dtFuef/8NDntvBvQ2kgVYNdIn9WsP3VXzqoXW1nWdaF+jzYZBsS43qV9JS5DFvi
27Tw56UTST3rNBPXX3OHKn/HWP27WUbEybYuWlV8Xdy/ZaKe2YIy/QG1y8NaumSeC6XfNTSdz1NL
jsiJSSbQuLxhBDQHkGzSgjWwJXBEK/ElngtymDmQ0z+CX9No+4PAeIB/bdAwCeD/Gh28K6qC+LwM
IsJtdBcchFJWnmM4N+YRKwSAVYLygRekhLhXZoCg8PSFCL3C6IEn40ZJMLNGHP3Nu6hQNdfIUxA4
YbriA0QfUNUpD1qi8GpxkHu+ULp2s/xxUVOxUJAU/cDgGcCKwaJPGY0djgFb4WvAy6r86mNRNRl4
Ykwa7220roJvM/hwu39QroHKz508GRMCsV5UZDItoKpAu7ul+5A/QojwRCpGYa0RWcNQcummGSq0
SujT9KJXGStsshF2kFNGnco3bl9/XIep8woazJDJmWESjPSToajuIXM3plNZx+np8Ln/ON/yXm5A
N6LZjOli204en1xuqzY3n8HqfXwQkmY7TdFzfQj5zE4OL+TS7zgK99Mwg1t/3rXM7gNTBJtiijtZ
wLH4lqmKN06XcVNeHPdZiT+agtS35YgYzCwdrnMobkpIYKIWhMy7Wr4PinDVGKTA/INScHJGHtiT
ABuoWJH1rX1RwZb6QKM0R3zSGSJDP5IjzuzxyIz/MAp2eLXKumOvid+t/vJOWmUqj2N9aGYFvVT9
PlNLelxXzsRRz0CWW74whQDBMnKDNsKvdCaG5oh3ayTZFQHm53M79rm1ZRBj1YmNpuaGbkeyXXf8
ouq9is4Apx9qGlK192YxR9wiKTiiLKrOZsYLyKxyfsP58Dn3mdHqsH8G+L7HeUkYK/40Ih2iJ8mh
Bbedjp1p2dv0QNPSmjRNatIj7FZIurk3Kl77zQqg+OLja0HZ0KhW+DYLpcqwaO4VTEvJKnK2wClo
pAfLfBUGJCInZAu5LMMuDKmbsTII5/lUPKk62CuPUx2a0CPjW2KcobllIt4vRdM7y3L9P4Xen9KT
xF+iHBnhW9d6OyRvThH57L6D/WcCgoH8WlNKHrTBYrx4BxWLJQ3skVTl4nL5o0hO5mxu28vZFPA0
0Xc5xK0gtyhoTWBO9t0BcDUqKSg/+RCjMETOKJLV51qa5xf95H66gcZLR81/o4cLifU5U6Dy0IQ9
luI9tPJUf1KGYUSWmlg9w+BDxyi09OTYV/jwkd97FKGNGIQXNyT2atk4hDvBi/wsE1eepl9nXN2J
+N30PX6hML6UD5rQ8i67Uyni63SEcXukrzcm05LO2ZTFA4E+iCjm4Iv0q9GD77GQPFWYVRuMLOf+
IRPUn1AnG8ik8TDNXju3A/LPMLg1Qbma8LvDvPYDyjbQ8ZqiuGhOVKtNwEbmf764QJ4fh29VBi4I
rS27URk3vU4aNa4r7+SGgYR+3ub1JJblWR1mL06OpAAQFT6dNwWjGwfUygVZ5nLmft6p5oPZL72s
0Zdasa8JXbeucJe9ljpk8UkBUHLQDS79uSqps3s6mTdTC720hYAeztyazJmirxLvI0CWIHjvGQO2
QZNcui/0KPLrI87404VokLrPhgbBVbRtQ0sQqkhxjCVRGcsguuKAKjRHVNvbmD+hTmc1TdW7zZfK
1erOLeGZ7dGf8tNvlVIRnl5fHigypQxd7yLJEYspxzqaHxzkj7U82OTino6TbP98EaK9tgX0vVxE
IOGdtYvwyhuCq9zedT8/cUWDfG1Xdh6fCMs9QT1odDCZngMHD4k7Tb+DottlZ6zZ9zY5IgpCH9RA
ye65Qo3/vbVoOYizdIL3nFsDXoG38ww81AJThewvvPeEwfGfVlnJLv477nKlyW9df/n/GpWRE0wl
kKuKoJGRfSxbXgrF4nAnAqHoADaKTR2jCSSMRks0FCbvTkTF5P408UmTH5hx0dRrjhC3a59LXie5
xWRSKK9Jk87wMA9vwRMUs66zO+7unYQ2hooDF9ATtaVWbpsCFFUnknCwu+jMCAwxaqFgchGe1Kvo
ub6xBf9qUKA4728kFzocDucFSQzb+PAluDVdU348+Cfb/L0bOTx5CBx7aSVEGqGodGyGgSwuoOgL
WEOBU+ldhWS+jwo/ppW0uF4to5wDz5M29PvHhzvT9jGl45B1rDMlY2d6xHLytlXk1xXf8zxKcnIr
8M06ZcHEGmKgH/SY2ZugbFS5U6mD29EO65Jfc5Yd/84tj8/SWlJ8o/9y2w58wK/UrPkwOOu+Kd0f
smfhqhc2/vU7UNZhg0uXi++KX0KDQ3JX86F/9vVvxQe3kyecLAN2tSj5Bo6knth6oGjFgeiqgKEW
on1/PYa7lbBiuyDkcDDMF/yLf/IEeETdIumdaR4+pqqP0jYW+e1su/09GyEwwoyz6XPp6qYp0gUZ
a+dcgCGwfQSZb6RzhbpEBj6tS+2q6YgCGvxGfPsU2QOYdNFCYNjh6+INxlWgDVfMrEucAQBUqGXp
BoqHU8RRm6nG6ciPBvpTLUpCpUmQ/bcOiHo/f4GiIiZTtH1ZMjdVdzv4sJ7nS2nZzhnxup3n6H2k
wAGkseEL5dtEpD9ksd1EZZ5e4MW1g/lzv38FOgbUb69UUpxTx0j/w9UAy5RD7Ts+/4eGEf96Vb25
PRDaZj+yQdX12tKh5fBpfRs8OshPwcta3PemDlOvjTrA58JTj9Tlu8uRBlplQKDF//a+f6k8nBL4
CavW7YEDAmCm8uf8Qq/dZBbI70qt+vLfnbMbqkaL2l6v18AzYTRM8YRO7j3xZPM74fCvpepXA1ND
JvEI18UprY5YDtEO6xzyDzgPuwTlBg2ihHO7/i5mkJ14pBa4I/5AznVgpuigxjpEFmqWVM1UQW16
PLfaB53FDO9HENw1ikHTjbOW9BPJoIkeT4lEMHZK5LivMWUGBxidF8TnoRZ04Yg50oGju65vFaKK
tRNcVMAv5I5ykhggPHdwIBlvyjkOfJBB+4HFyiDE6jkCj6Pv4UVY/5APye6v4zjFiIu9O3yKiRRQ
/7Cp/zcrHXIo0nvzeEdeykckdXM1rGCEEgg4Q3JcZNgfwt90JDgZu7dVoV7lzUHnwNP5G9uMTQkZ
MpPh7JJVylX9BsUdbgNtxeZjaDtk2scwkwvwm7LGecaADgaB5bIThnAtWJ/vZ3Z9U66J27fDFlJI
R2CUbvRqVoGwkfF7Av2dSzeMRKFjK9xUxDufdAe27abTxZrXTrpnIlIY8J2rgYSm2h9acxhiTrsm
2w5IRYu7K2xQ9w+/60qJ4DDpqx17js80QMXlcBJ5AFCWxmX75rp5rQmdPopk7FKGUwjDk4Af533T
LOIt/eoTT2qIlPvVIfDpgrti2dl3Rz/MTUwFAfJBETNk79twYex7afMJpDeE5KV4cpnvoZ0vfspB
PrQ+2vXZGAijboRIGB9avdXFDpN3ZI6vaH5sckkPaRzNZ4RxavUgzREb9aHf3xREYAJW1qT6Oz+K
5rvprwlmU9anF+QADcL1/Bb6vF8yxeaqLwlTtpb4w+/anyIqzvkbe6Gl5o065DOsczQxvqGDqaj/
PX96mixX4rq6NXC/eVrnaQjumzjHiYgOaDsa+dZYRy1YDKbdinZ4c48iiUYx4NxRy5PEuNgw7z7P
iEB+phchMkebkdS1x2NlEfkeX6vgebbO6KRATuz813zSt2FxzH/PKjBJdwnVRmq8C63p4ortUc3O
CVTi8hHACyiHpEU54UCsO5mpH+42zvqSIT4ikFCpE5X3x4h8Ef8Duw6Z0UgRxQRaBrFwNmkkOQrx
aaByTG8PH33udkp8tSj6Fkw1P9yqtQqdKB3MBEOQi7gTObszfnNv2exGxxRJ+EvhfRvpsbyfhf4L
5i1oSG+dsZJ5lznfaQa8GPo55w9hx10E77A6VMi//5MzOqfxBSLj8V+XiGY/caowVNlttL+RT2aq
mluXI+7CNxr40UrTCRq+ad9SiLCbXrQS4GpSwOIbxv98KkYYQeYGknZE35GuuOZZy1uTgmsSdA24
NOeebJJNVHeoq+sI94iADWoaJMESD+MavN9s21LLU1fpy9GLSEfgE2qgOIhnHiJZ8CdM5NVrhPXH
f/+COFBnsr9VzkT60EvoLBMgIVJotUvs5q0jUPhdvaTVQyfc8kE/1v61WWRci/kIQaSPsuR8LN/7
QFyhsSuHQxdg5fwCyj4nfnKPOHIlBomPbuMDEb3e62XQQCeoCiU1XZT8U29B3RKZLqRBk7QxteMY
a8Pg/I6D7ma2MLuBdK2Lt9P9hK7O34pAh+eGYxfljuWAWHPW0sqiQv1TSXaW/gXf674en2iE8HvZ
QqVo2Sqas5xbOR8tVuM9cWRJ0QAWiZzz1HPC8HgzA4QHh53/ML5QrXpdzMWYXeXK6LOu04ri0eyW
lxUeMVEQMdgfSaaNwyBDmaHZh3YnPJafeP+nPtRRcqqYgPjktESKNXcu0Q7ZbBBUaeVLm6XZp3rU
aoGehnLSnXC17UtFXKBD1pK9cKBu26DtOUkj2UDwsPzYqfnNPa3gf/LC2JR09Zq5bqr71Ya/mU8h
11PjbmG2m8Dh/zjrya827oSwuyYZQM6UBZU0p7U6N7/fXPo90bTVlQEj9k2hC/NF8EBNEA5lUpOz
KIbY0RjtoFvFc/YNzyCzIXcEKjXRpj/7ublPNn953Dy89oc0UftCJ/4ZRmt3FcFQQjLgwArJF/zB
VvzterOCPH1eFqQ6iDY2hWppZ4K3AJOYjMqL2UqfbfIKlUziXbDyOQ0q+1pad45IwCzoBPeF2ryd
fdy4QPkRKGqJ4C/b1LqPtLxLlAzynea2sUrRsBbeWdUwAAFTzZ8jYp/jlN+Y+JfKqP6shjgsFoFM
879bBLcUAtIElnyQyWOuWTSKm3lxBTxGa9PNaLJSWIXesmizoxuqA/J6DoB86k6jghG3lsQkw9Sy
EJgesahY/HWWkVgVkniehuqle9g6EkDYGEysRoxnboojn0FtX4e2jcTXZyatZ7pRZGyTPUw8CKcx
+/zRRA11Gw/EN1biZUtBDblizNkEl3lI8Q8g5kaV6YWo8bxnpJ543lQ0rulAx1TKQM40lsVY/+aM
QUJg1i0q3lDoqKoXYmiXsrxWQdXs43R6bXE0ppMhE0KSxsHr0dkyI1gGwwaa4XmYNDJNAcsdZYjg
kmS5QoJ2peGnWKIYY1bgNKoMIjom8qIIcIOPVEFPm3XpYuTY4/PUUZAOFhOT+1e+S2dCJwUvvnvU
sa6zmGSpabNN6c12rKyXCAi1gCKn4G0LXoEvVV1P1dpQkbtLuU2yl+iRvWFhGpdyjnn0xLQlH/Qd
hFXINEAjV7vuNs/zMo4N6sjvK7XXpotLvP4RyU1nJ9yRoD5j4nJ7peEk2++7DlSErQJsdGqAg3eI
btYcA7Bc/+dj01r+CcYsWLVnX1gLhG41qXXWMnkgCt7nB/Qo+ckIboQ3YVFO5tdlkB+Sn7sEAJXv
sKcyvXRMWQVhcbUVZnuFA1wl3vujNoKRapLVKrr9rB1mMbnOv2kKbUoZ65mm3hbLbUwITmxrZcWY
6Y4n4XZgFGDrAB0vQX0pToQ/jH3uaDGtnqVdpBcDAmsi5mv/mNcey0kYELBeEHCXgevv+uWQ4WfD
kZAgl8LbVebQGvBEC8xSaXkJfBLcJFsJbIJETgX6ags4bkBWCd1XF+3/C/jfAeFtn3aF/ATSka3C
pbSWlgF11ZQFS4NLUGQEA1LDhvvArI2kzYdgBkzUpvDj3vZ5v/4ChCXL/2F0QucQddXfqfpaQt4W
A0D3fkpoe9dvxR2XF+lgGERObYyj7jzHE/UBL7t/g0ntyeXqn7itpZfpeQ66vcMpnhtk+vUNHyWp
p3K9XiGMcxs1J75W6lS3x7TIHNyQn61+xY8Oc7yJskOw3SelHd9wwgQXFmztItL/PdxPuJ3t9Gjr
WIgjFttiqQ+8w0Bbd3uiBpfDCofyrjvTaM5YCVHCQMUfk3j5WYcG4EvVw7JmiBC70nCM6uPAnSQC
M6Fqg7cv+t/BIIQzCasbcN7cQ1jL9cc8IRniXwaWJP8jcgXP13uMKD4rqJN/rQdFmAXVjwhuwq5W
2iNd02F/54UW2k/6Z4+dwuDaq2iHXPjHwQ6+O+oqb8WbcdjVIEidk9iGoOsb6Ns7NqsQmH8llYgY
x0L3WNPOTVPQIGw/vtFR3F7z9AHr8xp/3XXNhLwdDweRxZIsQDsLQsctgnD4dkHXIyc2aPp5qTzh
5lyHpH/bBO746EG26zBoG7WAszWBvdMJNZn4+Bwf3bJVxCHUOoaJdfaEsGvOBkpdcYYzdi0L35tM
rlZReOAZR4mOT8CvdQ59ym545u2VZOEs116KHzn9XMpkAM+J+S/gj/fD0i5i3jvzFGUN8Z7twbAY
iymfFZjQ9gINGkIXkJHIVDmP25yYI3VV17zPjCK4AhU2ESPfs2sMvAa0ukP7abHZZVdTpgHRXC5b
hOSbJ39jqZsgc5QJt3CMTeFDwteG9z7LeLMRg77QAlXyV89vulzKTMQHzj9XbF21Rcl2hBQoTISX
qBGvfK9mnpcNAq04yfG4Cx9ic3dcvmlde1jv8D8qB5WF
`protect end_protected
